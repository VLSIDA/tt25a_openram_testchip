magic
tech sky130A
magscale 1 2
timestamp 1756238385
<< viali >>
rect 6193 44489 6227 44523
rect 6745 44489 6779 44523
rect 7297 44489 7331 44523
rect 7849 44489 7883 44523
rect 8401 44489 8435 44523
rect 8953 44489 8987 44523
rect 9505 44489 9539 44523
rect 10057 44489 10091 44523
rect 10517 44489 10551 44523
rect 10793 44489 10827 44523
rect 11161 44489 11195 44523
rect 11437 44489 11471 44523
rect 11713 44489 11747 44523
rect 12541 44489 12575 44523
rect 12817 44489 12851 44523
rect 20085 44489 20119 44523
rect 32413 44489 32447 44523
rect 11989 44421 12023 44455
rect 14381 44421 14415 44455
rect 27813 44421 27847 44455
rect 31217 44421 31251 44455
rect 46673 44421 46707 44455
rect 17049 44353 17083 44387
rect 17969 44353 18003 44387
rect 19809 44353 19843 44387
rect 22109 44353 22143 44387
rect 23949 44353 23983 44387
rect 24961 44353 24995 44387
rect 25697 44353 25731 44387
rect 27629 44353 27663 44387
rect 28641 44353 28675 44387
rect 29009 44353 29043 44387
rect 29837 44353 29871 44387
rect 30389 44353 30423 44387
rect 33885 44353 33919 44387
rect 36921 44353 36955 44387
rect 39405 44353 39439 44387
rect 42441 44353 42475 44387
rect 46305 44353 46339 44387
rect 12265 44285 12299 44319
rect 13277 44285 13311 44319
rect 14565 44285 14599 44319
rect 15117 44285 15151 44319
rect 15393 44285 15427 44319
rect 17141 44285 17175 44319
rect 18521 44285 18555 44319
rect 19625 44285 19659 44319
rect 20545 44285 20579 44319
rect 22937 44285 22971 44319
rect 23121 44285 23155 44319
rect 24133 44285 24167 44319
rect 27077 44285 27111 44319
rect 27997 44285 28031 44319
rect 31033 44285 31067 44319
rect 31401 44285 31435 44319
rect 31861 44285 31895 44319
rect 32045 44285 32079 44319
rect 32229 44285 32263 44319
rect 32597 44285 32631 44319
rect 34713 44285 34747 44319
rect 35541 44285 35575 44319
rect 38117 44285 38151 44319
rect 38577 44285 38611 44319
rect 38853 44285 38887 44319
rect 40509 44285 40543 44319
rect 41061 44285 41095 44319
rect 43361 44285 43395 44319
rect 44097 44285 44131 44319
rect 44465 44285 44499 44319
rect 46213 44285 46247 44319
rect 46857 44285 46891 44319
rect 14013 44217 14047 44251
rect 18705 44217 18739 44251
rect 19073 44217 19107 44251
rect 21097 44217 21131 44251
rect 21925 44217 21959 44251
rect 22661 44217 22695 44251
rect 25421 44217 25455 44251
rect 26893 44217 26927 44251
rect 28457 44217 28491 44251
rect 30481 44217 30515 44251
rect 33609 44217 33643 44251
rect 34161 44217 34195 44251
rect 36093 44217 36127 44251
rect 37105 44217 37139 44251
rect 37565 44217 37599 44251
rect 39681 44217 39715 44251
rect 41337 44217 41371 44251
rect 42257 44217 42291 44251
rect 43453 44217 43487 44251
rect 44741 44217 44775 44251
rect 47409 44217 47443 44251
rect 13185 44149 13219 44183
rect 13737 44149 13771 44183
rect 15025 44149 15059 44183
rect 15945 44149 15979 44183
rect 16405 44149 16439 44183
rect 17785 44149 17819 44183
rect 19257 44149 19291 44183
rect 19717 44149 19751 44183
rect 21557 44149 21591 44183
rect 22017 44149 22051 44183
rect 23673 44149 23707 44183
rect 24317 44149 24351 44183
rect 24685 44149 24719 44183
rect 24777 44149 24811 44183
rect 25329 44149 25363 44183
rect 26249 44149 26283 44183
rect 28089 44149 28123 44183
rect 28549 44149 28583 44183
rect 29653 44149 29687 44183
rect 31677 44149 31711 44183
rect 33241 44149 33275 44183
rect 33701 44149 33735 44183
rect 34989 44149 35023 44183
rect 35817 44149 35851 44183
rect 37013 44149 37047 44183
rect 37473 44149 37507 44183
rect 39957 44149 39991 44183
rect 40969 44149 41003 44183
rect 41429 44149 41463 44183
rect 41889 44149 41923 44183
rect 42349 44149 42383 44183
rect 42717 44149 42751 44183
rect 45753 44149 45787 44183
rect 46121 44149 46155 44183
rect 47133 44149 47167 44183
rect 14013 43945 14047 43979
rect 16865 43945 16899 43979
rect 16957 43945 16991 43979
rect 17325 43945 17359 43979
rect 17693 43945 17727 43979
rect 17785 43945 17819 43979
rect 18337 43945 18371 43979
rect 21741 43945 21775 43979
rect 23949 43945 23983 43979
rect 33425 43945 33459 43979
rect 36553 43945 36587 43979
rect 36737 43945 36771 43979
rect 39497 43945 39531 43979
rect 41429 43945 41463 43979
rect 46857 43945 46891 43979
rect 47409 43945 47443 43979
rect 11529 43877 11563 43911
rect 12909 43877 12943 43911
rect 13461 43877 13495 43911
rect 14105 43877 14139 43911
rect 14933 43877 14967 43911
rect 20821 43877 20855 43911
rect 22109 43877 22143 43911
rect 22201 43877 22235 43911
rect 24317 43877 24351 43911
rect 26157 43877 26191 43911
rect 27629 43877 27663 43911
rect 36093 43877 36127 43911
rect 36185 43877 36219 43911
rect 38209 43877 38243 43911
rect 41521 43877 41555 43911
rect 42165 43877 42199 43911
rect 44465 43877 44499 43911
rect 11437 43809 11471 43843
rect 11897 43809 11931 43843
rect 12817 43809 12851 43843
rect 13093 43809 13127 43843
rect 14841 43809 14875 43843
rect 15301 43809 15335 43843
rect 15853 43809 15887 43843
rect 16221 43809 16255 43843
rect 18521 43809 18555 43843
rect 18705 43809 18739 43843
rect 21649 43809 21683 43843
rect 27353 43809 27387 43843
rect 31677 43809 31711 43843
rect 35449 43809 35483 43843
rect 39129 43809 39163 43843
rect 44097 43809 44131 43843
rect 47869 43809 47903 43843
rect 52561 43809 52595 43843
rect 52745 43809 52779 43843
rect 53941 43809 53975 43843
rect 11621 43741 11655 43775
rect 12449 43741 12483 43775
rect 14197 43741 14231 43775
rect 15025 43741 15059 43775
rect 17141 43741 17175 43775
rect 17877 43741 17911 43775
rect 19257 43741 19291 43775
rect 21097 43741 21131 43775
rect 22385 43741 22419 43775
rect 23121 43741 23155 43775
rect 23397 43741 23431 43775
rect 24041 43741 24075 43775
rect 26433 43741 26467 43775
rect 27077 43741 27111 43775
rect 29193 43741 29227 43775
rect 29469 43741 29503 43775
rect 31217 43741 31251 43775
rect 31953 43741 31987 43775
rect 33517 43741 33551 43775
rect 33793 43741 33827 43775
rect 35909 43741 35943 43775
rect 38485 43741 38519 43775
rect 40969 43741 41003 43775
rect 41245 43741 41279 43775
rect 41889 43741 41923 43775
rect 44281 43741 44315 43775
rect 45109 43741 45143 43775
rect 45385 43741 45419 43775
rect 47501 43741 47535 43775
rect 47685 43741 47719 43775
rect 13277 43673 13311 43707
rect 21465 43673 21499 43707
rect 43637 43673 43671 43707
rect 52929 43673 52963 43707
rect 11069 43605 11103 43639
rect 13645 43605 13679 43639
rect 14473 43605 14507 43639
rect 16497 43605 16531 43639
rect 19349 43605 19383 43639
rect 22569 43605 22603 43639
rect 25789 43605 25823 43639
rect 26065 43605 26099 43639
rect 29101 43605 29135 43639
rect 35265 43605 35299 43639
rect 35541 43605 35575 43639
rect 38577 43605 38611 43639
rect 43821 43605 43855 43639
rect 47041 43605 47075 43639
rect 48513 43605 48547 43639
rect 52285 43605 52319 43639
rect 53665 43605 53699 43639
rect 17417 43401 17451 43435
rect 17509 43401 17543 43435
rect 20453 43401 20487 43435
rect 22569 43401 22603 43435
rect 25605 43401 25639 43435
rect 28825 43401 28859 43435
rect 29561 43401 29595 43435
rect 34161 43401 34195 43435
rect 34989 43401 35023 43435
rect 36369 43401 36403 43435
rect 40785 43401 40819 43435
rect 43545 43401 43579 43435
rect 48789 43401 48823 43435
rect 53941 43401 53975 43435
rect 25697 43333 25731 43367
rect 29285 43333 29319 43367
rect 43453 43333 43487 43367
rect 15117 43265 15151 43299
rect 15669 43265 15703 43299
rect 18429 43265 18463 43299
rect 20821 43265 20855 43299
rect 23857 43265 23891 43299
rect 26341 43265 26375 43299
rect 26801 43265 26835 43299
rect 27813 43265 27847 43299
rect 28273 43265 28307 43299
rect 30113 43265 30147 43299
rect 31769 43265 31803 43299
rect 34805 43265 34839 43299
rect 35541 43265 35575 43299
rect 38761 43265 38795 43299
rect 40509 43265 40543 43299
rect 41429 43265 41463 43299
rect 41705 43265 41739 43299
rect 44005 43265 44039 43299
rect 44097 43265 44131 43299
rect 45385 43265 45419 43299
rect 46857 43265 46891 43299
rect 47317 43265 47351 43299
rect 50629 43265 50663 43299
rect 52377 43265 52411 43299
rect 53021 43265 53055 43299
rect 10701 43197 10735 43231
rect 15393 43197 15427 43231
rect 18153 43197 18187 43231
rect 18705 43197 18739 43231
rect 22661 43197 22695 43231
rect 23673 43197 23707 43231
rect 26985 43197 27019 43231
rect 28365 43197 28399 43231
rect 28457 43197 28491 43231
rect 29929 43197 29963 43231
rect 31309 43197 31343 43231
rect 33885 43197 33919 43231
rect 34529 43197 34563 43231
rect 35357 43197 35391 43231
rect 38117 43197 38151 43231
rect 38577 43197 38611 43231
rect 40325 43197 40359 43231
rect 41153 43197 41187 43231
rect 45109 43197 45143 43231
rect 47041 43197 47075 43231
rect 53297 43197 53331 43231
rect 53849 43197 53883 43231
rect 10977 43129 11011 43163
rect 15945 43129 15979 43163
rect 18981 43129 19015 43163
rect 21097 43129 21131 43163
rect 24133 43129 24167 43163
rect 26893 43129 26927 43163
rect 27537 43129 27571 43163
rect 29101 43129 29135 43163
rect 30481 43129 30515 43163
rect 32045 43129 32079 43163
rect 33701 43129 33735 43163
rect 35449 43129 35483 43163
rect 37841 43129 37875 43163
rect 39405 43129 39439 43163
rect 41981 43129 42015 43163
rect 43913 43129 43947 43163
rect 50905 43129 50939 43163
rect 12449 43061 12483 43095
rect 13645 43061 13679 43095
rect 17785 43061 17819 43095
rect 18245 43061 18279 43095
rect 22845 43061 22879 43095
rect 23029 43061 23063 43095
rect 26065 43061 26099 43095
rect 26157 43061 26191 43095
rect 27353 43061 27387 43095
rect 30021 43061 30055 43095
rect 30573 43061 30607 43095
rect 31401 43061 31435 43095
rect 33517 43061 33551 43095
rect 34621 43061 34655 43095
rect 38209 43061 38243 43095
rect 38669 43061 38703 43095
rect 39497 43061 39531 43095
rect 39957 43061 39991 43095
rect 40417 43061 40451 43095
rect 41245 43061 41279 43095
rect 52469 43061 52503 43095
rect 53389 43061 53423 43095
rect 11345 42857 11379 42891
rect 11713 42857 11747 42891
rect 14565 42857 14599 42891
rect 15209 42857 15243 42891
rect 16865 42857 16899 42891
rect 19349 42857 19383 42891
rect 20085 42857 20119 42891
rect 20453 42857 20487 42891
rect 20545 42857 20579 42891
rect 21925 42857 21959 42891
rect 25789 42857 25823 42891
rect 25881 42857 25915 42891
rect 26249 42857 26283 42891
rect 26433 42857 26467 42891
rect 27169 42857 27203 42891
rect 27997 42857 28031 42891
rect 29929 42857 29963 42891
rect 32689 42857 32723 42891
rect 33057 42857 33091 42891
rect 34345 42857 34379 42891
rect 34805 42857 34839 42891
rect 36093 42857 36127 42891
rect 39497 42857 39531 42891
rect 40141 42857 40175 42891
rect 40509 42857 40543 42891
rect 41705 42857 41739 42891
rect 44097 42857 44131 42891
rect 46765 42857 46799 42891
rect 47869 42857 47903 42891
rect 48237 42857 48271 42891
rect 51273 42857 51307 42891
rect 51641 42857 51675 42891
rect 15577 42789 15611 42823
rect 15669 42789 15703 42823
rect 17877 42789 17911 42823
rect 19901 42789 19935 42823
rect 22385 42789 22419 42823
rect 23121 42789 23155 42823
rect 27077 42789 27111 42823
rect 29101 42789 29135 42823
rect 30297 42789 30331 42823
rect 36185 42789 36219 42823
rect 37013 42789 37047 42823
rect 41337 42789 41371 42823
rect 11805 42721 11839 42755
rect 15117 42721 15151 42755
rect 16129 42721 16163 42755
rect 17325 42721 17359 42755
rect 17601 42721 17635 42755
rect 22293 42721 22327 42755
rect 25053 42721 25087 42755
rect 26617 42721 26651 42755
rect 27905 42721 27939 42755
rect 28365 42721 28399 42755
rect 30389 42721 30423 42755
rect 32229 42721 32263 42755
rect 33517 42721 33551 42755
rect 34437 42721 34471 42755
rect 37105 42721 37139 42755
rect 39589 42721 39623 42755
rect 47317 42721 47351 42755
rect 47409 42721 47443 42755
rect 48697 42721 48731 42755
rect 9505 42653 9539 42687
rect 11989 42653 12023 42687
rect 12817 42653 12851 42687
rect 13093 42653 13127 42687
rect 15761 42653 15795 42687
rect 16957 42653 16991 42687
rect 17141 42653 17175 42687
rect 20637 42653 20671 42687
rect 21373 42653 21407 42687
rect 22109 42653 22143 42687
rect 22845 42653 22879 42687
rect 24593 42653 24627 42687
rect 25145 42653 25179 42687
rect 25329 42653 25363 42687
rect 25697 42653 25731 42687
rect 27261 42653 27295 42687
rect 28089 42653 28123 42687
rect 28917 42653 28951 42687
rect 29653 42653 29687 42687
rect 30481 42653 30515 42687
rect 31677 42653 31711 42687
rect 32505 42653 32539 42687
rect 32597 42653 32631 42687
rect 33609 42653 33643 42687
rect 33701 42653 33735 42687
rect 34253 42653 34287 42687
rect 35909 42653 35943 42687
rect 36829 42653 36863 42687
rect 37565 42653 37599 42687
rect 38853 42653 38887 42687
rect 39681 42653 39715 42687
rect 40601 42653 40635 42687
rect 40785 42653 40819 42687
rect 41061 42653 41095 42687
rect 41245 42653 41279 42687
rect 41889 42653 41923 42687
rect 42165 42653 42199 42687
rect 44189 42653 44223 42687
rect 44281 42653 44315 42687
rect 45017 42653 45051 42687
rect 45293 42653 45327 42687
rect 47133 42653 47167 42687
rect 48329 42653 48363 42687
rect 48421 42653 48455 42687
rect 49249 42653 49283 42687
rect 51733 42653 51767 42687
rect 51917 42653 51951 42687
rect 52193 42653 52227 42687
rect 52469 42653 52503 42687
rect 54217 42653 54251 42687
rect 33149 42585 33183 42619
rect 36553 42585 36587 42619
rect 38301 42585 38335 42619
rect 43729 42585 43763 42619
rect 47777 42585 47811 42619
rect 8953 42517 8987 42551
rect 16313 42517 16347 42551
rect 16497 42517 16531 42551
rect 22753 42517 22787 42551
rect 24685 42517 24719 42551
rect 26709 42517 26743 42551
rect 27537 42517 27571 42551
rect 37473 42517 37507 42551
rect 38209 42517 38243 42551
rect 39129 42517 39163 42551
rect 43637 42517 43671 42551
rect 11713 42313 11747 42347
rect 12541 42313 12575 42347
rect 17601 42313 17635 42347
rect 19809 42313 19843 42347
rect 20177 42313 20211 42347
rect 24777 42313 24811 42347
rect 25605 42313 25639 42347
rect 28365 42313 28399 42347
rect 32891 42313 32925 42347
rect 33241 42313 33275 42347
rect 34161 42313 34195 42347
rect 35909 42313 35943 42347
rect 41245 42313 41279 42347
rect 44465 42313 44499 42347
rect 45569 42313 45603 42347
rect 52009 42313 52043 42347
rect 52101 42313 52135 42347
rect 22109 42245 22143 42279
rect 53113 42245 53147 42279
rect 9965 42177 9999 42211
rect 13001 42177 13035 42211
rect 13185 42177 13219 42211
rect 15393 42177 15427 42211
rect 15669 42177 15703 42211
rect 18061 42177 18095 42211
rect 18153 42177 18187 42211
rect 19165 42177 19199 42211
rect 22017 42177 22051 42211
rect 22569 42177 22603 42211
rect 22661 42177 22695 42211
rect 23581 42177 23615 42211
rect 24133 42177 24167 42211
rect 26157 42177 26191 42211
rect 26249 42177 26283 42211
rect 26617 42177 26651 42211
rect 33149 42177 33183 42211
rect 33793 42177 33827 42211
rect 34713 42177 34747 42211
rect 38301 42177 38335 42211
rect 38393 42177 38427 42211
rect 39313 42177 39347 42211
rect 45017 42177 45051 42211
rect 46121 42177 46155 42211
rect 48237 42177 48271 42211
rect 48421 42177 48455 42211
rect 50169 42177 50203 42211
rect 50997 42177 51031 42211
rect 51457 42177 51491 42211
rect 52653 42177 52687 42211
rect 9689 42109 9723 42143
rect 13737 42109 13771 42143
rect 14565 42109 14599 42143
rect 19441 42109 19475 42143
rect 22477 42109 22511 42143
rect 23305 42109 23339 42143
rect 23397 42109 23431 42143
rect 24317 42109 24351 42143
rect 26065 42109 26099 42143
rect 29377 42109 29411 42143
rect 33609 42109 33643 42143
rect 35081 42109 35115 42143
rect 37749 42109 37783 42143
rect 38209 42109 38243 42143
rect 44925 42109 44959 42143
rect 46489 42109 46523 42143
rect 49985 42109 50019 42143
rect 52469 42109 52503 42143
rect 53389 42109 53423 42143
rect 10241 42041 10275 42075
rect 11989 42041 12023 42075
rect 12357 42041 12391 42075
rect 12909 42041 12943 42075
rect 17509 42041 17543 42075
rect 17969 42041 18003 42075
rect 21741 42041 21775 42075
rect 26893 42041 26927 42075
rect 37473 42041 37507 42075
rect 39589 42041 39623 42075
rect 41521 42041 41555 42075
rect 41889 42041 41923 42075
rect 43637 42041 43671 42075
rect 44833 42041 44867 42075
rect 45293 42041 45327 42075
rect 45937 42041 45971 42075
rect 46765 42041 46799 42075
rect 50077 42041 50111 42075
rect 50813 42041 50847 42075
rect 53665 42041 53699 42075
rect 54033 42041 54067 42075
rect 55781 42041 55815 42075
rect 9045 41973 9079 42007
rect 14381 41973 14415 42007
rect 15117 41973 15151 42007
rect 17141 41973 17175 42007
rect 19349 41973 19383 42007
rect 20269 41973 20303 42007
rect 22937 41973 22971 42007
rect 24409 41973 24443 42007
rect 25697 41973 25731 42007
rect 29101 41973 29135 42007
rect 31401 41973 31435 42007
rect 33701 41973 33735 42007
rect 36001 41973 36035 42007
rect 37841 41973 37875 42007
rect 41061 41973 41095 42007
rect 46029 41973 46063 42007
rect 49065 41973 49099 42007
rect 49617 41973 49651 42007
rect 50445 41973 50479 42007
rect 50905 41973 50939 42007
rect 51549 41973 51583 42007
rect 51641 41973 51675 42007
rect 52561 41973 52595 42007
rect 56057 41973 56091 42007
rect 9505 41769 9539 41803
rect 9965 41769 9999 41803
rect 15577 41769 15611 41803
rect 15669 41769 15703 41803
rect 17785 41769 17819 41803
rect 22017 41769 22051 41803
rect 22477 41769 22511 41803
rect 24777 41769 24811 41803
rect 25237 41769 25271 41803
rect 25605 41769 25639 41803
rect 28181 41769 28215 41803
rect 33241 41769 33275 41803
rect 33701 41769 33735 41803
rect 36277 41769 36311 41803
rect 36737 41769 36771 41803
rect 37197 41769 37231 41803
rect 41889 41769 41923 41803
rect 42349 41769 42383 41803
rect 43177 41769 43211 41803
rect 43545 41769 43579 41803
rect 45753 41769 45787 41803
rect 47593 41769 47627 41803
rect 48053 41769 48087 41803
rect 48145 41769 48179 41803
rect 48513 41769 48547 41803
rect 53021 41769 53055 41803
rect 17049 41701 17083 41735
rect 18245 41701 18279 41735
rect 20177 41701 20211 41735
rect 22569 41701 22603 41735
rect 23305 41701 23339 41735
rect 25697 41701 25731 41735
rect 26709 41701 26743 41735
rect 34529 41701 34563 41735
rect 38853 41701 38887 41735
rect 40509 41701 40543 41735
rect 43085 41701 43119 41735
rect 44189 41701 44223 41735
rect 46121 41701 46155 41735
rect 48605 41701 48639 41735
rect 49709 41701 49743 41735
rect 7757 41633 7791 41667
rect 10057 41633 10091 41667
rect 17141 41633 17175 41667
rect 17693 41633 17727 41667
rect 18153 41633 18187 41667
rect 19533 41633 19567 41667
rect 21557 41633 21591 41667
rect 21649 41633 21683 41667
rect 26433 41633 26467 41667
rect 28641 41633 28675 41667
rect 29101 41633 29135 41667
rect 33333 41633 33367 41667
rect 35725 41633 35759 41667
rect 36185 41633 36219 41667
rect 37105 41633 37139 41667
rect 37565 41633 37599 41667
rect 38577 41633 38611 41667
rect 42257 41633 42291 41667
rect 44097 41633 44131 41667
rect 45109 41633 45143 41667
rect 47685 41633 47719 41667
rect 52561 41633 52595 41667
rect 53757 41633 53791 41667
rect 55229 41633 55263 41667
rect 55965 41633 55999 41667
rect 8033 41565 8067 41599
rect 10241 41565 10275 41599
rect 11529 41565 11563 41599
rect 11805 41565 11839 41599
rect 13277 41565 13311 41599
rect 13921 41565 13955 41599
rect 14565 41565 14599 41599
rect 15853 41565 15887 41599
rect 16865 41565 16899 41599
rect 18337 41565 18371 41599
rect 19165 41565 19199 41599
rect 21465 41565 21499 41599
rect 22661 41565 22695 41599
rect 23029 41565 23063 41599
rect 25789 41565 25823 41599
rect 28733 41565 28767 41599
rect 28825 41565 28859 41599
rect 29745 41565 29779 41599
rect 33057 41565 33091 41599
rect 34069 41565 34103 41599
rect 35173 41565 35207 41599
rect 36369 41565 36403 41599
rect 37289 41565 37323 41599
rect 37841 41565 37875 41599
rect 40325 41565 40359 41599
rect 42533 41565 42567 41599
rect 43361 41565 43395 41599
rect 44373 41565 44407 41599
rect 46213 41565 46247 41599
rect 46397 41565 46431 41599
rect 47409 41565 47443 41599
rect 48697 41565 48731 41599
rect 49433 41565 49467 41599
rect 51457 41565 51491 41599
rect 52653 41565 52687 41599
rect 52837 41565 52871 41599
rect 53665 41565 53699 41599
rect 54309 41565 54343 41599
rect 55321 41565 55355 41599
rect 55505 41565 55539 41599
rect 56609 41565 56643 41599
rect 9597 41497 9631 41531
rect 15117 41497 15151 41531
rect 28273 41497 28307 41531
rect 44557 41497 44591 41531
rect 13369 41429 13403 41463
rect 15209 41429 15243 41463
rect 17509 41429 17543 41463
rect 18613 41429 18647 41463
rect 20085 41429 20119 41463
rect 22109 41429 22143 41463
rect 35817 41429 35851 41463
rect 38485 41429 38519 41463
rect 42717 41429 42751 41463
rect 43729 41429 43763 41463
rect 52193 41429 52227 41463
rect 54861 41429 54895 41463
rect 10149 41225 10183 41259
rect 11805 41225 11839 41259
rect 16773 41225 16807 41259
rect 29009 41225 29043 41259
rect 32965 41225 32999 41259
rect 51365 41225 51399 41259
rect 56517 41225 56551 41259
rect 20177 41157 20211 41191
rect 23489 41157 23523 41191
rect 36645 41157 36679 41191
rect 44465 41157 44499 41191
rect 46213 41157 46247 41191
rect 7665 41089 7699 41123
rect 8401 41089 8435 41123
rect 10885 41089 10919 41123
rect 12357 41089 12391 41123
rect 13185 41089 13219 41123
rect 14105 41089 14139 41123
rect 17877 41089 17911 41123
rect 18061 41089 18095 41123
rect 19257 41089 19291 41123
rect 24501 41089 24535 41123
rect 26617 41089 26651 41123
rect 29653 41089 29687 41123
rect 33793 41089 33827 41123
rect 34897 41089 34931 41123
rect 36737 41089 36771 41123
rect 37933 41089 37967 41123
rect 38669 41089 38703 41123
rect 39773 41089 39807 41123
rect 39957 41089 39991 41123
rect 42441 41089 42475 41123
rect 44189 41089 44223 41123
rect 45109 41089 45143 41123
rect 46029 41089 46063 41123
rect 53849 41089 53883 41123
rect 10609 41021 10643 41055
rect 12173 41021 12207 41055
rect 13001 41021 13035 41055
rect 13093 41021 13127 41055
rect 15025 41021 15059 41055
rect 17325 41021 17359 41055
rect 17785 41021 17819 41055
rect 19073 41021 19107 41055
rect 21741 41021 21775 41055
rect 24225 41021 24259 41055
rect 28273 41021 28307 41055
rect 29377 41021 29411 41055
rect 30481 41021 30515 41055
rect 31861 41021 31895 41055
rect 32321 41021 32355 41055
rect 34713 41021 34747 41055
rect 37749 41021 37783 41055
rect 42257 41021 42291 41055
rect 44833 41021 44867 41055
rect 46765 41021 46799 41055
rect 46949 41021 46983 41055
rect 49617 41021 49651 41055
rect 51457 41021 51491 41055
rect 54769 41021 54803 41055
rect 56977 41021 57011 41055
rect 57161 41021 57195 41055
rect 57253 41021 57287 41055
rect 57437 41021 57471 41055
rect 7849 40953 7883 40987
rect 8677 40953 8711 40987
rect 12265 40953 12299 40987
rect 14013 40953 14047 40987
rect 15301 40953 15335 40987
rect 19165 40953 19199 40987
rect 21649 40953 21683 40987
rect 22017 40953 22051 40987
rect 24685 40953 24719 40987
rect 32873 40953 32907 40987
rect 33517 40953 33551 40987
rect 35173 40953 35207 40987
rect 40509 40953 40543 40987
rect 42717 40953 42751 40987
rect 44925 40953 44959 40987
rect 47225 40953 47259 40987
rect 49893 40953 49927 40987
rect 53205 40953 53239 40987
rect 55045 40953 55079 40987
rect 56609 40953 56643 40987
rect 7757 40885 7791 40919
rect 8217 40885 8251 40919
rect 10241 40885 10275 40919
rect 10701 40885 10735 40919
rect 12633 40885 12667 40919
rect 13553 40885 13587 40919
rect 13921 40885 13955 40919
rect 17417 40885 17451 40919
rect 18705 40885 18739 40919
rect 23857 40885 23891 40919
rect 24317 40885 24351 40919
rect 26157 40885 26191 40919
rect 29469 40885 29503 40919
rect 29837 40885 29871 40919
rect 31309 40885 31343 40919
rect 33149 40885 33183 40919
rect 33609 40885 33643 40919
rect 34161 40885 34195 40919
rect 37289 40885 37323 40919
rect 37657 40885 37691 40919
rect 38117 40885 38151 40919
rect 38485 40885 38519 40919
rect 38577 40885 38611 40919
rect 39313 40885 39347 40919
rect 39681 40885 39715 40919
rect 45385 40885 45419 40919
rect 45753 40885 45787 40919
rect 45845 40885 45879 40919
rect 48697 40885 48731 40919
rect 53297 40885 53331 40919
rect 53665 40885 53699 40919
rect 53757 40885 53791 40919
rect 7941 40681 7975 40715
rect 8309 40681 8343 40715
rect 11345 40681 11379 40715
rect 15209 40681 15243 40715
rect 15577 40681 15611 40715
rect 15669 40681 15703 40715
rect 22017 40681 22051 40715
rect 22937 40681 22971 40715
rect 29469 40681 29503 40715
rect 29929 40681 29963 40715
rect 31033 40681 31067 40715
rect 33517 40681 33551 40715
rect 33977 40681 34011 40715
rect 37197 40681 37231 40715
rect 41061 40681 41095 40715
rect 42073 40681 42107 40715
rect 9045 40613 9079 40647
rect 12449 40613 12483 40647
rect 23213 40613 23247 40647
rect 23765 40613 23799 40647
rect 25697 40613 25731 40647
rect 34805 40613 34839 40647
rect 38485 40613 38519 40647
rect 39497 40613 39531 40647
rect 42625 40613 42659 40647
rect 45109 40613 45143 40647
rect 47777 40613 47811 40647
rect 50261 40613 50295 40647
rect 52469 40613 52503 40647
rect 10793 40545 10827 40579
rect 11437 40545 11471 40579
rect 14565 40545 14599 40579
rect 16129 40545 16163 40579
rect 18061 40545 18095 40579
rect 18521 40545 18555 40579
rect 21649 40545 21683 40579
rect 23489 40545 23523 40579
rect 25789 40545 25823 40579
rect 26433 40545 26467 40579
rect 27353 40545 27387 40579
rect 27629 40545 27663 40579
rect 29837 40545 29871 40579
rect 31769 40545 31803 40579
rect 39221 40545 39255 40579
rect 41981 40545 42015 40579
rect 47869 40545 47903 40579
rect 48973 40545 49007 40579
rect 49801 40545 49835 40579
rect 52193 40545 52227 40579
rect 8401 40477 8435 40511
rect 8585 40477 8619 40511
rect 8769 40477 8803 40511
rect 11529 40477 11563 40511
rect 12173 40477 12207 40511
rect 14197 40477 14231 40511
rect 15761 40477 15795 40511
rect 16405 40477 16439 40511
rect 18613 40477 18647 40511
rect 18797 40477 18831 40511
rect 20729 40477 20763 40511
rect 21005 40477 21039 40511
rect 21465 40477 21499 40511
rect 21557 40477 21591 40511
rect 22109 40477 22143 40511
rect 25237 40477 25271 40511
rect 25973 40477 26007 40511
rect 27077 40477 27111 40511
rect 27905 40477 27939 40511
rect 30113 40477 30147 40511
rect 31125 40477 31159 40511
rect 31309 40477 31343 40511
rect 32045 40477 32079 40511
rect 34069 40477 34103 40511
rect 34161 40477 34195 40511
rect 41613 40477 41647 40511
rect 42349 40477 42383 40511
rect 44833 40477 44867 40511
rect 48053 40477 48087 40511
rect 49065 40477 49099 40511
rect 49157 40477 49191 40511
rect 49525 40477 49559 40511
rect 49709 40477 49743 40511
rect 53941 40477 53975 40511
rect 54585 40477 54619 40511
rect 54861 40477 54895 40511
rect 56609 40477 56643 40511
rect 18153 40409 18187 40443
rect 33609 40409 33643 40443
rect 36093 40409 36127 40443
rect 47409 40409 47443 40443
rect 50169 40409 50203 40443
rect 51549 40409 51583 40443
rect 10977 40341 11011 40375
rect 15117 40341 15151 40375
rect 17877 40341 17911 40375
rect 19257 40341 19291 40375
rect 22753 40341 22787 40375
rect 25329 40341 25363 40375
rect 29377 40341 29411 40375
rect 30665 40341 30699 40375
rect 40969 40341 41003 40375
rect 44097 40341 44131 40375
rect 46581 40341 46615 40375
rect 48605 40341 48639 40375
rect 15227 40137 15261 40171
rect 17067 40137 17101 40171
rect 19336 40137 19370 40171
rect 20913 40137 20947 40171
rect 21833 40137 21867 40171
rect 24856 40137 24890 40171
rect 27064 40137 27098 40171
rect 28549 40137 28583 40171
rect 30008 40137 30042 40171
rect 31493 40137 31527 40171
rect 33069 40137 33103 40171
rect 34161 40137 34195 40171
rect 35344 40137 35378 40171
rect 37644 40137 37678 40171
rect 39129 40137 39163 40171
rect 43269 40137 43303 40171
rect 46581 40137 46615 40171
rect 47948 40137 47982 40171
rect 55597 40137 55631 40171
rect 9321 40001 9355 40035
rect 9505 40001 9539 40035
rect 9781 40001 9815 40035
rect 11529 40001 11563 40035
rect 13737 40001 13771 40035
rect 15577 40001 15611 40035
rect 18245 40001 18279 40035
rect 21557 40001 21591 40035
rect 22293 40001 22327 40035
rect 22477 40001 22511 40035
rect 22661 40001 22695 40035
rect 23305 40001 23339 40035
rect 24593 40001 24627 40035
rect 34713 40001 34747 40035
rect 36829 40001 36863 40035
rect 37381 40001 37415 40035
rect 42257 40001 42291 40035
rect 43085 40001 43119 40035
rect 43913 40001 43947 40035
rect 44833 40001 44867 40035
rect 45109 40001 45143 40035
rect 47225 40001 47259 40035
rect 47685 40001 47719 40035
rect 49709 40001 49743 40035
rect 53849 40001 53883 40035
rect 54125 40001 54159 40035
rect 54861 40001 54895 40035
rect 56241 40001 56275 40035
rect 7665 39933 7699 39967
rect 12817 39933 12851 39967
rect 15485 39933 15519 39967
rect 17325 39933 17359 39967
rect 19073 39933 19107 39967
rect 21281 39933 21315 39967
rect 24409 39933 24443 39967
rect 26801 39933 26835 39967
rect 29745 39933 29779 39967
rect 33333 39933 33367 39967
rect 35081 39933 35115 39967
rect 39773 39933 39807 39967
rect 41981 39933 42015 39967
rect 55045 39933 55079 39967
rect 55965 39933 55999 39967
rect 8217 39865 8251 39899
rect 9045 39865 9079 39899
rect 13369 39865 13403 39899
rect 22201 39865 22235 39899
rect 34529 39865 34563 39899
rect 40049 39865 40083 39899
rect 50721 39865 50755 39899
rect 52101 39865 52135 39899
rect 56057 39865 56091 39899
rect 8677 39797 8711 39831
rect 9137 39797 9171 39831
rect 17601 39797 17635 39831
rect 17969 39797 18003 39831
rect 18061 39797 18095 39831
rect 20821 39797 20855 39831
rect 21373 39797 21407 39831
rect 23857 39797 23891 39831
rect 26341 39797 26375 39831
rect 31585 39797 31619 39831
rect 34621 39797 34655 39831
rect 41521 39797 41555 39831
rect 41613 39797 41647 39831
rect 42073 39797 42107 39831
rect 43637 39797 43671 39831
rect 43729 39797 43763 39831
rect 46673 39797 46707 39831
rect 49433 39797 49467 39831
rect 49893 39797 49927 39831
rect 49985 39797 50019 39831
rect 50353 39797 50387 39831
rect 55137 39797 55171 39831
rect 55505 39797 55539 39831
rect 18429 39593 18463 39627
rect 20453 39593 20487 39627
rect 21281 39593 21315 39627
rect 22109 39593 22143 39627
rect 22477 39593 22511 39627
rect 24041 39593 24075 39627
rect 25145 39593 25179 39627
rect 25513 39593 25547 39627
rect 28457 39593 28491 39627
rect 28825 39593 28859 39627
rect 31033 39593 31067 39627
rect 33425 39593 33459 39627
rect 33885 39593 33919 39627
rect 36093 39593 36127 39627
rect 36553 39593 36587 39627
rect 38577 39593 38611 39627
rect 38945 39593 38979 39627
rect 42901 39593 42935 39627
rect 43729 39593 43763 39627
rect 44189 39593 44223 39627
rect 46121 39593 46155 39627
rect 46489 39593 46523 39627
rect 52377 39593 52411 39627
rect 8861 39525 8895 39559
rect 9689 39525 9723 39559
rect 11437 39525 11471 39559
rect 15577 39525 15611 39559
rect 16957 39525 16991 39559
rect 19165 39525 19199 39559
rect 36185 39525 36219 39559
rect 37013 39525 37047 39559
rect 39037 39525 39071 39559
rect 41429 39525 41463 39559
rect 43269 39525 43303 39559
rect 50261 39525 50295 39559
rect 50629 39525 50663 39559
rect 51365 39525 51399 39559
rect 52837 39525 52871 39559
rect 9137 39457 9171 39491
rect 9597 39457 9631 39491
rect 11345 39457 11379 39491
rect 13737 39457 13771 39491
rect 14197 39457 14231 39491
rect 14289 39457 14323 39491
rect 16681 39457 16715 39491
rect 21649 39457 21683 39491
rect 21741 39457 21775 39491
rect 29837 39457 29871 39491
rect 31585 39457 31619 39491
rect 33793 39457 33827 39491
rect 36737 39457 36771 39491
rect 41705 39457 41739 39491
rect 42441 39457 42475 39491
rect 42533 39457 42567 39491
rect 44097 39457 44131 39491
rect 45661 39457 45695 39491
rect 47041 39457 47075 39491
rect 51181 39457 51215 39491
rect 52745 39457 52779 39491
rect 55873 39457 55907 39491
rect 56425 39457 56459 39491
rect 58541 39457 58575 39491
rect 7389 39389 7423 39423
rect 9781 39389 9815 39423
rect 11621 39389 11655 39423
rect 13461 39389 13495 39423
rect 14381 39389 14415 39423
rect 15301 39389 15335 39423
rect 15485 39389 15519 39423
rect 21833 39389 21867 39423
rect 22569 39389 22603 39423
rect 22661 39389 22695 39423
rect 23857 39389 23891 39423
rect 23949 39389 23983 39423
rect 25605 39389 25639 39423
rect 25789 39389 25823 39423
rect 26985 39389 27019 39423
rect 27721 39389 27755 39423
rect 28917 39389 28951 39423
rect 29009 39389 29043 39423
rect 30757 39389 30791 39423
rect 30941 39389 30975 39423
rect 31861 39389 31895 39423
rect 33977 39389 34011 39423
rect 35909 39389 35943 39423
rect 39129 39389 39163 39423
rect 42625 39389 42659 39423
rect 43361 39389 43395 39423
rect 43453 39389 43487 39423
rect 44281 39389 44315 39423
rect 45109 39389 45143 39423
rect 45477 39389 45511 39423
rect 45569 39389 45603 39423
rect 46581 39389 46615 39423
rect 46765 39389 46799 39423
rect 48513 39389 48547 39423
rect 50537 39389 50571 39423
rect 53021 39389 53055 39423
rect 53849 39389 53883 39423
rect 55965 39389 55999 39423
rect 56149 39389 56183 39423
rect 56977 39389 57011 39423
rect 58817 39389 58851 39423
rect 60933 39389 60967 39423
rect 10977 39321 11011 39355
rect 13829 39321 13863 39355
rect 15945 39321 15979 39355
rect 31401 39321 31435 39355
rect 39957 39321 39991 39355
rect 46029 39321 46063 39355
rect 9229 39253 9263 39287
rect 11989 39253 12023 39287
rect 24409 39253 24443 39287
rect 26433 39253 26467 39287
rect 27169 39253 27203 39287
rect 29285 39253 29319 39287
rect 33333 39253 33367 39287
rect 38485 39253 38519 39287
rect 42073 39253 42107 39287
rect 47685 39253 47719 39287
rect 53205 39253 53239 39287
rect 55505 39253 55539 39287
rect 60289 39253 60323 39287
rect 60381 39253 60415 39287
rect 21189 39049 21223 39083
rect 23673 39049 23707 39083
rect 43361 39049 43395 39083
rect 45293 39049 45327 39083
rect 46121 39049 46155 39083
rect 48697 39049 48731 39083
rect 15301 38981 15335 39015
rect 21097 38981 21131 39015
rect 25605 38981 25639 39015
rect 31585 38981 31619 39015
rect 37657 38981 37691 39015
rect 39313 38981 39347 39015
rect 58909 38981 58943 39015
rect 8493 38913 8527 38947
rect 10517 38913 10551 38947
rect 10609 38913 10643 38947
rect 12817 38913 12851 38947
rect 12909 38913 12943 38947
rect 13553 38913 13587 38947
rect 16773 38913 16807 38947
rect 19349 38913 19383 38947
rect 21925 38913 21959 38947
rect 23857 38913 23891 38947
rect 24133 38913 24167 38947
rect 26341 38913 26375 38947
rect 27629 38913 27663 38947
rect 28549 38913 28583 38947
rect 30205 38913 30239 38947
rect 30941 38913 30975 38947
rect 32229 38913 32263 38947
rect 35633 38913 35667 38947
rect 38209 38913 38243 38947
rect 39865 38913 39899 38947
rect 40601 38913 40635 38947
rect 40693 38913 40727 38947
rect 41521 38913 41555 38947
rect 43269 38913 43303 38947
rect 43913 38913 43947 38947
rect 45017 38913 45051 38947
rect 49157 38913 49191 38947
rect 49249 38913 49283 38947
rect 50445 38913 50479 38947
rect 53941 38913 53975 38947
rect 55045 38913 55079 38947
rect 58633 38913 58667 38947
rect 59461 38913 59495 38947
rect 60473 38913 60507 38947
rect 8217 38845 8251 38879
rect 13001 38845 13035 38879
rect 16037 38845 16071 38879
rect 21741 38845 21775 38879
rect 26065 38845 26099 38879
rect 30757 38845 30791 38879
rect 32045 38845 32079 38879
rect 32413 38845 32447 38879
rect 32965 38845 32999 38879
rect 33977 38845 34011 38879
rect 34161 38845 34195 38879
rect 35541 38845 35575 38879
rect 38117 38845 38151 38879
rect 38485 38845 38519 38879
rect 39681 38845 39715 38879
rect 45845 38845 45879 38879
rect 47869 38845 47903 38879
rect 49065 38845 49099 38879
rect 51457 38845 51491 38879
rect 58541 38845 58575 38879
rect 59277 38845 59311 38879
rect 8769 38777 8803 38811
rect 10885 38777 10919 38811
rect 13829 38777 13863 38811
rect 18521 38777 18555 38811
rect 19625 38777 19659 38811
rect 22201 38777 22235 38811
rect 27445 38777 27479 38811
rect 30849 38777 30883 38811
rect 31953 38777 31987 38811
rect 33333 38777 33367 38811
rect 35909 38777 35943 38811
rect 37473 38777 37507 38811
rect 38025 38777 38059 38811
rect 41797 38777 41831 38811
rect 44833 38777 44867 38811
rect 47593 38777 47627 38811
rect 50261 38777 50295 38811
rect 50905 38777 50939 38811
rect 53665 38777 53699 38811
rect 55321 38777 55355 38811
rect 58449 38777 58483 38811
rect 59921 38777 59955 38811
rect 7573 38709 7607 38743
rect 12357 38709 12391 38743
rect 13369 38709 13403 38743
rect 15485 38709 15519 38743
rect 25697 38709 25731 38743
rect 26157 38709 26191 38743
rect 27077 38709 27111 38743
rect 27537 38709 27571 38743
rect 27905 38709 27939 38743
rect 28273 38709 28307 38743
rect 28365 38709 28399 38743
rect 29561 38709 29595 38743
rect 29929 38709 29963 38743
rect 30021 38709 30055 38743
rect 30389 38709 30423 38743
rect 34805 38709 34839 38743
rect 34897 38709 34931 38743
rect 37381 38709 37415 38743
rect 39129 38709 39163 38743
rect 39773 38709 39807 38743
rect 40141 38709 40175 38743
rect 40509 38709 40543 38743
rect 44465 38709 44499 38743
rect 44925 38709 44959 38743
rect 49893 38709 49927 38743
rect 50353 38709 50387 38743
rect 52193 38709 52227 38743
rect 56793 38709 56827 38743
rect 58081 38709 58115 38743
rect 59369 38709 59403 38743
rect 8861 38505 8895 38539
rect 9229 38505 9263 38539
rect 9597 38505 9631 38539
rect 10793 38505 10827 38539
rect 14013 38505 14047 38539
rect 14473 38505 14507 38539
rect 15669 38505 15703 38539
rect 20177 38505 20211 38539
rect 20545 38505 20579 38539
rect 21649 38505 21683 38539
rect 23121 38505 23155 38539
rect 23489 38505 23523 38539
rect 30757 38505 30791 38539
rect 35357 38505 35391 38539
rect 35449 38505 35483 38539
rect 35817 38505 35851 38539
rect 36737 38505 36771 38539
rect 37105 38505 37139 38539
rect 38209 38505 38243 38539
rect 40417 38505 40451 38539
rect 40877 38505 40911 38539
rect 45661 38505 45695 38539
rect 47409 38505 47443 38539
rect 47777 38505 47811 38539
rect 48421 38505 48455 38539
rect 48789 38505 48823 38539
rect 48881 38505 48915 38539
rect 53297 38505 53331 38539
rect 53665 38505 53699 38539
rect 60289 38505 60323 38539
rect 10425 38437 10459 38471
rect 11989 38437 12023 38471
rect 14105 38437 14139 38471
rect 27353 38437 27387 38471
rect 29193 38437 29227 38471
rect 36277 38437 36311 38471
rect 43453 38437 43487 38471
rect 44097 38437 44131 38471
rect 49893 38437 49927 38471
rect 54493 38437 54527 38471
rect 59553 38437 59587 38471
rect 7113 38369 7147 38403
rect 11529 38369 11563 38403
rect 12541 38369 12575 38403
rect 15577 38369 15611 38403
rect 16497 38369 16531 38403
rect 17601 38369 17635 38403
rect 22477 38369 22511 38403
rect 24133 38369 24167 38403
rect 28917 38369 28951 38403
rect 34897 38369 34931 38403
rect 36185 38369 36219 38403
rect 37197 38369 37231 38403
rect 40785 38369 40819 38403
rect 43821 38369 43855 38403
rect 49617 38369 49651 38403
rect 54401 38369 54435 38403
rect 55137 38369 55171 38403
rect 57437 38369 57471 38403
rect 7389 38301 7423 38335
rect 9689 38301 9723 38335
rect 9873 38301 9907 38335
rect 10241 38301 10275 38335
rect 10333 38301 10367 38335
rect 11621 38301 11655 38335
rect 11805 38301 11839 38335
rect 13921 38301 13955 38335
rect 15853 38301 15887 38335
rect 16589 38301 16623 38335
rect 16681 38301 16715 38335
rect 19901 38301 19935 38335
rect 20085 38301 20119 38335
rect 21741 38301 21775 38335
rect 21925 38301 21959 38335
rect 23581 38301 23615 38335
rect 23765 38301 23799 38335
rect 24409 38301 24443 38335
rect 27077 38301 27111 38335
rect 30665 38301 30699 38335
rect 31309 38301 31343 38335
rect 34621 38301 34655 38335
rect 35541 38301 35575 38335
rect 36369 38301 36403 38335
rect 37289 38301 37323 38335
rect 39681 38301 39715 38335
rect 39957 38301 39991 38335
rect 41061 38301 41095 38335
rect 43729 38301 43763 38335
rect 45569 38301 45603 38335
rect 46213 38301 46247 38335
rect 47133 38301 47167 38335
rect 47317 38301 47351 38335
rect 48973 38301 49007 38335
rect 52745 38301 52779 38335
rect 53021 38301 53055 38335
rect 53205 38301 53239 38335
rect 54677 38301 54711 38335
rect 56885 38301 56919 38335
rect 57161 38301 57195 38335
rect 57805 38301 57839 38335
rect 59829 38301 59863 38335
rect 60381 38301 60415 38335
rect 60565 38301 60599 38335
rect 22201 38233 22235 38267
rect 34989 38233 35023 38267
rect 52193 38233 52227 38267
rect 54033 38233 54067 38267
rect 11161 38165 11195 38199
rect 15209 38165 15243 38199
rect 16129 38165 16163 38199
rect 21281 38165 21315 38199
rect 25881 38165 25915 38199
rect 28825 38165 28859 38199
rect 33149 38165 33183 38199
rect 41981 38165 42015 38199
rect 51365 38165 51399 38199
rect 53849 38165 53883 38199
rect 59921 38165 59955 38199
rect 7481 37961 7515 37995
rect 17233 37961 17267 37995
rect 18705 37961 18739 37995
rect 19809 37961 19843 37995
rect 23857 37961 23891 37995
rect 33793 37961 33827 37995
rect 36921 37961 36955 37995
rect 41245 37961 41279 37995
rect 42809 37961 42843 37995
rect 43637 37961 43671 37995
rect 44557 37961 44591 37995
rect 51825 37961 51859 37995
rect 57805 37961 57839 37995
rect 60657 37961 60691 37995
rect 16681 37893 16715 37927
rect 28273 37893 28307 37927
rect 29009 37893 29043 37927
rect 35081 37893 35115 37927
rect 56057 37893 56091 37927
rect 56885 37893 56919 37927
rect 8125 37825 8159 37859
rect 8401 37825 8435 37859
rect 10425 37825 10459 37859
rect 10701 37825 10735 37859
rect 10977 37825 11011 37859
rect 14565 37825 14599 37859
rect 14657 37825 14691 37859
rect 14933 37825 14967 37859
rect 15209 37825 15243 37859
rect 19349 37825 19383 37859
rect 20453 37825 20487 37859
rect 20637 37825 20671 37859
rect 24501 37825 24535 37859
rect 26525 37825 26559 37859
rect 26801 37825 26835 37859
rect 29929 37825 29963 37859
rect 32034 37825 32068 37859
rect 34253 37825 34287 37859
rect 34437 37825 34471 37859
rect 38209 37825 38243 37859
rect 38577 37825 38611 37859
rect 39957 37825 39991 37859
rect 40785 37825 40819 37859
rect 42257 37825 42291 37859
rect 43085 37825 43119 37859
rect 48421 37825 48455 37859
rect 50077 37825 50111 37859
rect 54585 37825 54619 37859
rect 55505 37825 55539 37859
rect 56241 37825 56275 37859
rect 57253 37825 57287 37859
rect 58173 37825 58207 37859
rect 60105 37825 60139 37859
rect 7849 37757 7883 37791
rect 18521 37757 18555 37791
rect 20177 37757 20211 37791
rect 24685 37757 24719 37791
rect 29561 37757 29595 37791
rect 34529 37757 34563 37791
rect 35633 37757 35667 37791
rect 38669 37757 38703 37791
rect 39681 37757 39715 37791
rect 39773 37757 39807 37791
rect 40509 37757 40543 37791
rect 41797 37757 41831 37791
rect 42441 37757 42475 37791
rect 43177 37757 43211 37791
rect 43269 37757 43303 37791
rect 46305 37757 46339 37791
rect 48690 37757 48724 37791
rect 49341 37757 49375 37791
rect 55689 37757 55723 37791
rect 57897 37757 57931 37791
rect 60289 37757 60323 37791
rect 63417 37757 63451 37791
rect 8677 37689 8711 37723
rect 12725 37689 12759 37723
rect 20913 37689 20947 37723
rect 24961 37689 24995 37723
rect 30205 37689 30239 37723
rect 32321 37689 32355 37723
rect 35357 37689 35391 37723
rect 38761 37689 38795 37723
rect 40601 37689 40635 37723
rect 46029 37689 46063 37723
rect 50353 37689 50387 37723
rect 52561 37689 52595 37723
rect 54309 37689 54343 37723
rect 56425 37689 56459 37723
rect 56517 37689 56551 37723
rect 57437 37689 57471 37723
rect 7941 37621 7975 37655
rect 14105 37621 14139 37655
rect 14473 37621 14507 37655
rect 19073 37621 19107 37655
rect 19165 37621 19199 37655
rect 20269 37621 20303 37655
rect 22385 37621 22419 37655
rect 24225 37621 24259 37655
rect 24317 37621 24351 37655
rect 26433 37621 26467 37655
rect 31677 37621 31711 37655
rect 34897 37621 34931 37655
rect 39129 37621 39163 37655
rect 39313 37621 39347 37655
rect 40141 37621 40175 37655
rect 42349 37621 42383 37655
rect 46949 37621 46983 37655
rect 48789 37621 48823 37655
rect 55597 37621 55631 37655
rect 57345 37621 57379 37655
rect 59645 37621 59679 37655
rect 60197 37621 60231 37655
rect 64061 37621 64095 37655
rect 9045 37417 9079 37451
rect 9505 37417 9539 37451
rect 10977 37417 11011 37451
rect 12265 37417 12299 37451
rect 12725 37417 12759 37451
rect 15301 37417 15335 37451
rect 19073 37417 19107 37451
rect 21373 37417 21407 37451
rect 21741 37417 21775 37451
rect 25513 37417 25547 37451
rect 25881 37417 25915 37451
rect 25973 37417 26007 37451
rect 26433 37417 26467 37451
rect 26893 37417 26927 37451
rect 27905 37417 27939 37451
rect 28273 37417 28307 37451
rect 30389 37417 30423 37451
rect 30757 37417 30791 37451
rect 32413 37417 32447 37451
rect 32873 37417 32907 37451
rect 33241 37417 33275 37451
rect 36553 37417 36587 37451
rect 44741 37417 44775 37451
rect 45201 37417 45235 37451
rect 45661 37417 45695 37451
rect 46029 37417 46063 37451
rect 47777 37417 47811 37451
rect 48237 37417 48271 37451
rect 48605 37417 48639 37451
rect 49985 37417 50019 37451
rect 50905 37417 50939 37451
rect 51273 37417 51307 37451
rect 51365 37417 51399 37451
rect 52193 37417 52227 37451
rect 52561 37417 52595 37451
rect 53205 37417 53239 37451
rect 53757 37417 53791 37451
rect 54125 37417 54159 37451
rect 56701 37417 56735 37451
rect 56793 37417 56827 37451
rect 62497 37417 62531 37451
rect 9413 37349 9447 37383
rect 12633 37349 12667 37383
rect 13829 37349 13863 37383
rect 32781 37349 32815 37383
rect 33701 37349 33735 37383
rect 35081 37349 35115 37383
rect 36737 37349 36771 37383
rect 40233 37349 40267 37383
rect 45569 37349 45603 37383
rect 47317 37349 47351 37383
rect 50445 37349 50479 37383
rect 52653 37349 52687 37383
rect 59645 37349 59679 37383
rect 11345 37281 11379 37315
rect 11437 37281 11471 37315
rect 13553 37281 13587 37315
rect 16773 37281 16807 37315
rect 19165 37281 19199 37315
rect 21833 37281 21867 37315
rect 26801 37281 26835 37315
rect 28365 37281 28399 37315
rect 30849 37281 30883 37315
rect 31585 37281 31619 37315
rect 32137 37281 32171 37315
rect 33609 37281 33643 37315
rect 34805 37281 34839 37315
rect 39957 37281 39991 37315
rect 44833 37281 44867 37315
rect 47409 37281 47443 37315
rect 49801 37281 49835 37315
rect 50353 37281 50387 37315
rect 56057 37281 56091 37315
rect 57621 37281 57655 37315
rect 64245 37281 64279 37315
rect 9597 37213 9631 37247
rect 11529 37213 11563 37247
rect 12817 37213 12851 37247
rect 17049 37213 17083 37247
rect 19257 37213 19291 37247
rect 21925 37213 21959 37247
rect 26157 37213 26191 37247
rect 27077 37213 27111 37247
rect 28549 37213 28583 37247
rect 31033 37213 31067 37247
rect 33057 37213 33091 37247
rect 33885 37213 33919 37247
rect 38485 37213 38519 37247
rect 44557 37213 44591 37247
rect 45477 37213 45511 37247
rect 47225 37213 47259 37247
rect 47961 37213 47995 37247
rect 48145 37213 48179 37247
rect 50537 37213 50571 37247
rect 51549 37213 51583 37247
rect 52837 37213 52871 37247
rect 53573 37213 53607 37247
rect 53665 37213 53699 37247
rect 56609 37213 56643 37247
rect 57897 37213 57931 37247
rect 63969 37213 64003 37247
rect 65993 37213 66027 37247
rect 18705 37145 18739 37179
rect 57161 37145 57195 37179
rect 18521 37077 18555 37111
rect 41705 37077 41739 37111
rect 65441 37077 65475 37111
rect 63877 36873 63911 36907
rect 64429 36737 64463 36771
rect 65257 36737 65291 36771
rect 64245 36669 64279 36703
rect 65073 36669 65107 36703
rect 64337 36601 64371 36635
rect 64705 36533 64739 36567
rect 65165 36533 65199 36567
rect 64153 36261 64187 36295
rect 63877 36125 63911 36159
rect 65625 35989 65659 36023
rect 65073 35785 65107 35819
rect 64797 35649 64831 35683
rect 65533 35649 65567 35683
rect 65625 35649 65659 35683
rect 64613 35581 64647 35615
rect 65441 35513 65475 35547
rect 64245 35445 64279 35479
rect 64705 35445 64739 35479
rect 64153 35173 64187 35207
rect 63877 35037 63911 35071
rect 65625 34901 65659 34935
rect 64705 34697 64739 34731
rect 64613 34629 64647 34663
rect 63969 34561 64003 34595
rect 65165 34561 65199 34595
rect 65257 34561 65291 34595
rect 64153 34493 64187 34527
rect 64245 34425 64279 34459
rect 65073 34425 65107 34459
rect 65165 34153 65199 34187
rect 65717 34017 65751 34051
rect 65165 33473 65199 33507
rect 65993 33473 66027 33507
rect 64889 33337 64923 33371
rect 65441 33337 65475 33371
rect 64521 33269 64555 33303
rect 64981 33269 65015 33303
rect 65809 33065 65843 33099
rect 64337 32997 64371 33031
rect 64061 32929 64095 32963
rect 65073 32521 65107 32555
rect 64521 32385 64555 32419
rect 64613 32385 64647 32419
rect 64705 32317 64739 32351
rect 64981 31977 65015 32011
rect 65349 31977 65383 32011
rect 64889 31841 64923 31875
rect 64797 31773 64831 31807
rect 65533 31773 65567 31807
rect 66085 31773 66119 31807
rect 65165 31433 65199 31467
rect 63877 31229 63911 31263
rect 65165 30889 65199 30923
rect 63877 30753 63911 30787
rect 64061 30209 64095 30243
rect 64337 30073 64371 30107
rect 65809 30005 65843 30039
rect 65349 29801 65383 29835
rect 65717 29801 65751 29835
rect 65809 29801 65843 29835
rect 64889 29733 64923 29767
rect 64981 29665 65015 29699
rect 65073 29597 65107 29631
rect 65901 29597 65935 29631
rect 64521 29461 64555 29495
rect 65809 29257 65843 29291
rect 64061 29121 64095 29155
rect 64337 29121 64371 29155
rect 64797 28713 64831 28747
rect 65165 28713 65199 28747
rect 64705 28645 64739 28679
rect 65441 28645 65475 28679
rect 65993 28577 66027 28611
rect 64613 28509 64647 28543
rect 64429 28169 64463 28203
rect 65073 27625 65107 27659
rect 64981 27489 65015 27523
rect 65257 27421 65291 27455
rect 64613 27285 64647 27319
rect 64061 26945 64095 26979
rect 64337 26809 64371 26843
rect 65809 26741 65843 26775
rect 64613 26537 64647 26571
rect 65073 26537 65107 26571
rect 64981 26401 65015 26435
rect 65441 26401 65475 26435
rect 65993 26401 66027 26435
rect 65257 26333 65291 26367
rect 63969 25313 64003 25347
rect 64981 25313 65015 25347
rect 65441 25313 65475 25347
rect 65073 25245 65107 25279
rect 65165 25245 65199 25279
rect 65993 25245 66027 25279
rect 64613 25109 64647 25143
rect 63877 24701 63911 24735
rect 65165 24565 65199 24599
rect 65165 24361 65199 24395
rect 63877 24293 63911 24327
rect 64061 23613 64095 23647
rect 64337 23545 64371 23579
rect 65809 23477 65843 23511
rect 65257 23273 65291 23307
rect 64797 23205 64831 23239
rect 64429 23137 64463 23171
rect 64889 23137 64923 23171
rect 64705 23069 64739 23103
rect 64613 22729 64647 22763
rect 64337 22525 64371 22559
rect 65349 22457 65383 22491
rect 65717 22457 65751 22491
rect 65809 22185 65843 22219
rect 64061 22049 64095 22083
rect 64337 21981 64371 22015
rect 65993 21437 66027 21471
rect 64981 21369 65015 21403
rect 65349 21369 65383 21403
rect 65441 21301 65475 21335
rect 64613 21097 64647 21131
rect 64981 21097 65015 21131
rect 65073 20893 65107 20927
rect 65257 20893 65291 20927
rect 65165 20417 65199 20451
rect 65073 20349 65107 20383
rect 64613 20213 64647 20247
rect 64981 20213 65015 20247
rect 64061 19805 64095 19839
rect 64337 19805 64371 19839
rect 65809 19669 65843 19703
rect 64613 19465 64647 19499
rect 65257 19329 65291 19363
rect 65073 19261 65107 19295
rect 65993 19261 66027 19295
rect 64981 19193 65015 19227
rect 65441 19193 65475 19227
rect 64981 18785 65015 18819
rect 65441 18785 65475 18819
rect 65073 18717 65107 18751
rect 65257 18717 65291 18751
rect 65993 18717 66027 18751
rect 64613 18581 64647 18615
rect 64337 18241 64371 18275
rect 64061 18173 64095 18207
rect 65809 18037 65843 18071
rect 64797 17833 64831 17867
rect 65349 17833 65383 17867
rect 65717 17833 65751 17867
rect 64889 17765 64923 17799
rect 65809 17697 65843 17731
rect 64705 17629 64739 17663
rect 65901 17629 65935 17663
rect 65257 17561 65291 17595
rect 64613 17289 64647 17323
rect 64981 16609 65015 16643
rect 65441 16609 65475 16643
rect 65993 16609 66027 16643
rect 65073 16541 65107 16575
rect 65165 16541 65199 16575
rect 64613 16405 64647 16439
rect 65809 16201 65843 16235
rect 64061 16065 64095 16099
rect 64337 16065 64371 16099
rect 64981 15657 65015 15691
rect 65349 15657 65383 15691
rect 64889 15589 64923 15623
rect 64797 15453 64831 15487
rect 64705 15113 64739 15147
rect 64061 12801 64095 12835
rect 64337 12801 64371 12835
rect 66085 12801 66119 12835
rect 65809 12393 65843 12427
rect 64061 12189 64095 12223
rect 64337 12189 64371 12223
rect 64521 11849 64555 11883
rect 65349 11849 65383 11883
rect 65165 11713 65199 11747
rect 65901 11713 65935 11747
rect 64981 11645 65015 11679
rect 65717 11577 65751 11611
rect 64889 11509 64923 11543
rect 65809 11509 65843 11543
rect 65441 11305 65475 11339
rect 65993 11169 66027 11203
rect 64613 10693 64647 10727
rect 65165 10625 65199 10659
rect 65073 10557 65107 10591
rect 64981 10421 65015 10455
rect 64061 10013 64095 10047
rect 64337 10013 64371 10047
rect 65809 9877 65843 9911
rect 65191 9537 65225 9571
rect 65993 9469 66027 9503
rect 65441 9401 65475 9435
rect 64889 9333 64923 9367
rect 64981 9333 65015 9367
rect 65349 9333 65383 9367
rect 64613 9129 64647 9163
rect 64981 9129 65015 9163
rect 65073 8925 65107 8959
rect 65257 8925 65291 8959
rect 65257 8449 65291 8483
rect 65073 8381 65107 8415
rect 65993 8381 66027 8415
rect 64981 8313 65015 8347
rect 65441 8313 65475 8347
rect 64613 8245 64647 8279
rect 64337 7973 64371 8007
rect 64061 7905 64095 7939
rect 65809 7701 65843 7735
rect 65257 7497 65291 7531
rect 64705 7361 64739 7395
rect 64797 7361 64831 7395
rect 64889 7293 64923 7327
rect 65993 7293 66027 7327
rect 65441 7157 65475 7191
rect 65257 6953 65291 6987
rect 63877 6817 63911 6851
rect 64521 6817 64555 6851
rect 64705 6817 64739 6851
rect 65349 6817 65383 6851
rect 64153 6749 64187 6783
rect 65533 6749 65567 6783
rect 64889 6613 64923 6647
rect 64705 6409 64739 6443
rect 64061 6273 64095 6307
rect 65257 6273 65291 6307
rect 64153 6205 64187 6239
rect 65073 6205 65107 6239
rect 65165 6205 65199 6239
rect 64245 6137 64279 6171
rect 64613 6069 64647 6103
rect 64337 5865 64371 5899
rect 64705 5865 64739 5899
rect 64245 5729 64279 5763
rect 64429 5661 64463 5695
rect 63877 5525 63911 5559
rect 65809 5321 65843 5355
rect 64061 5185 64095 5219
rect 64337 5185 64371 5219
rect 65625 4777 65659 4811
rect 63877 4641 63911 4675
rect 64153 4573 64187 4607
rect 64134 4233 64168 4267
rect 63877 4029 63911 4063
rect 65625 3893 65659 3927
rect 64153 3689 64187 3723
rect 64613 3689 64647 3723
rect 65165 3689 65199 3723
rect 64245 3621 64279 3655
rect 65073 3553 65107 3587
rect 64061 3485 64095 3519
rect 65349 3485 65383 3519
rect 64705 3349 64739 3383
rect 63877 3145 63911 3179
rect 64061 3009 64095 3043
rect 64337 2873 64371 2907
rect 65809 2805 65843 2839
rect 63877 2601 63911 2635
rect 64705 2601 64739 2635
rect 65165 2601 65199 2635
rect 64429 2465 64463 2499
rect 65257 2465 65291 2499
rect 65349 2397 65383 2431
rect 64797 2261 64831 2295
rect 65441 2057 65475 2091
rect 65349 1989 65383 2023
rect 64705 1921 64739 1955
rect 64889 1921 64923 1955
rect 65993 1853 66027 1887
rect 64981 1785 65015 1819
rect 64705 1513 64739 1547
rect 65257 1513 65291 1547
rect 65165 1377 65199 1411
rect 65441 1309 65475 1343
rect 64797 1241 64831 1275
rect 65441 969 65475 1003
rect 65993 833 66027 867
<< metal1 >>
rect 21266 44956 21272 45008
rect 21324 44996 21330 45008
rect 39390 44996 39396 45008
rect 21324 44968 39396 44996
rect 21324 44956 21330 44968
rect 39390 44956 39396 44968
rect 39448 44956 39454 45008
rect 15102 44752 15108 44804
rect 15160 44792 15166 44804
rect 22830 44792 22836 44804
rect 15160 44764 22836 44792
rect 15160 44752 15166 44764
rect 22830 44752 22836 44764
rect 22888 44752 22894 44804
rect 14550 44684 14556 44736
rect 14608 44724 14614 44736
rect 21450 44724 21456 44736
rect 14608 44696 21456 44724
rect 14608 44684 14614 44696
rect 21450 44684 21456 44696
rect 21508 44724 21514 44736
rect 22002 44724 22008 44736
rect 21508 44696 22008 44724
rect 21508 44684 21514 44696
rect 22002 44684 22008 44696
rect 22060 44684 22066 44736
rect 23290 44684 23296 44736
rect 23348 44724 23354 44736
rect 26418 44724 26424 44736
rect 23348 44696 26424 44724
rect 23348 44684 23354 44696
rect 26418 44684 26424 44696
rect 26476 44684 26482 44736
rect 29086 44684 29092 44736
rect 29144 44724 29150 44736
rect 32398 44724 32404 44736
rect 29144 44696 32404 44724
rect 29144 44684 29150 44696
rect 32398 44684 32404 44696
rect 32456 44684 32462 44736
rect 552 44634 66424 44656
rect 552 44582 1998 44634
rect 2050 44582 2062 44634
rect 2114 44582 2126 44634
rect 2178 44582 2190 44634
rect 2242 44582 2254 44634
rect 2306 44582 49998 44634
rect 50050 44582 50062 44634
rect 50114 44582 50126 44634
rect 50178 44582 50190 44634
rect 50242 44582 50254 44634
rect 50306 44582 66424 44634
rect 552 44560 66424 44582
rect 6178 44480 6184 44532
rect 6236 44480 6242 44532
rect 6730 44480 6736 44532
rect 6788 44480 6794 44532
rect 7282 44480 7288 44532
rect 7340 44480 7346 44532
rect 7834 44480 7840 44532
rect 7892 44480 7898 44532
rect 8386 44480 8392 44532
rect 8444 44480 8450 44532
rect 8938 44480 8944 44532
rect 8996 44480 9002 44532
rect 9490 44480 9496 44532
rect 9548 44480 9554 44532
rect 10042 44480 10048 44532
rect 10100 44480 10106 44532
rect 10502 44480 10508 44532
rect 10560 44480 10566 44532
rect 10778 44480 10784 44532
rect 10836 44480 10842 44532
rect 11146 44480 11152 44532
rect 11204 44480 11210 44532
rect 11422 44480 11428 44532
rect 11480 44480 11486 44532
rect 11698 44480 11704 44532
rect 11756 44480 11762 44532
rect 12526 44480 12532 44532
rect 12584 44480 12590 44532
rect 12805 44523 12863 44529
rect 12805 44489 12817 44523
rect 12851 44520 12863 44523
rect 15194 44520 15200 44532
rect 12851 44492 15200 44520
rect 12851 44489 12863 44492
rect 12805 44483 12863 44489
rect 15194 44480 15200 44492
rect 15252 44480 15258 44532
rect 18414 44480 18420 44532
rect 18472 44520 18478 44532
rect 18472 44492 19840 44520
rect 18472 44480 18478 44492
rect 11977 44455 12035 44461
rect 11977 44421 11989 44455
rect 12023 44452 12035 44455
rect 13814 44452 13820 44464
rect 12023 44424 13820 44452
rect 12023 44421 12035 44424
rect 11977 44415 12035 44421
rect 13814 44412 13820 44424
rect 13872 44412 13878 44464
rect 14369 44455 14427 44461
rect 14369 44421 14381 44455
rect 14415 44452 14427 44455
rect 16482 44452 16488 44464
rect 14415 44424 16488 44452
rect 14415 44421 14427 44424
rect 14369 44415 14427 44421
rect 16482 44412 16488 44424
rect 16540 44412 16546 44464
rect 19702 44452 19708 44464
rect 16960 44424 19708 44452
rect 16960 44384 16988 44424
rect 19702 44412 19708 44424
rect 19760 44412 19766 44464
rect 13280 44356 16988 44384
rect 17037 44387 17095 44393
rect 13280 44325 13308 44356
rect 17037 44353 17049 44387
rect 17083 44384 17095 44387
rect 17218 44384 17224 44396
rect 17083 44356 17224 44384
rect 17083 44353 17095 44356
rect 17037 44347 17095 44353
rect 17218 44344 17224 44356
rect 17276 44344 17282 44396
rect 17957 44387 18015 44393
rect 17957 44353 17969 44387
rect 18003 44384 18015 44387
rect 19518 44384 19524 44396
rect 18003 44356 19524 44384
rect 18003 44353 18015 44356
rect 17957 44347 18015 44353
rect 19518 44344 19524 44356
rect 19576 44344 19582 44396
rect 19812 44393 19840 44492
rect 20070 44480 20076 44532
rect 20128 44480 20134 44532
rect 26326 44520 26332 44532
rect 22940 44492 26332 44520
rect 19886 44412 19892 44464
rect 19944 44452 19950 44464
rect 21634 44452 21640 44464
rect 19944 44424 21640 44452
rect 19944 44412 19950 44424
rect 21634 44412 21640 44424
rect 21692 44452 21698 44464
rect 21692 44424 22232 44452
rect 21692 44412 21698 44424
rect 19797 44387 19855 44393
rect 19797 44353 19809 44387
rect 19843 44353 19855 44387
rect 21910 44384 21916 44396
rect 19797 44347 19855 44353
rect 19904 44356 21916 44384
rect 12253 44319 12311 44325
rect 12253 44285 12265 44319
rect 12299 44285 12311 44319
rect 12253 44279 12311 44285
rect 13265 44319 13323 44325
rect 13265 44285 13277 44319
rect 13311 44285 13323 44319
rect 14366 44316 14372 44328
rect 13265 44279 13323 44285
rect 13556 44288 14372 44316
rect 12268 44248 12296 44279
rect 13556 44248 13584 44288
rect 14366 44276 14372 44288
rect 14424 44276 14430 44328
rect 14550 44276 14556 44328
rect 14608 44276 14614 44328
rect 15102 44276 15108 44328
rect 15160 44276 15166 44328
rect 15378 44276 15384 44328
rect 15436 44276 15442 44328
rect 17129 44319 17187 44325
rect 17129 44285 17141 44319
rect 17175 44316 17187 44319
rect 17770 44316 17776 44328
rect 17175 44288 17776 44316
rect 17175 44285 17187 44288
rect 17129 44279 17187 44285
rect 17770 44276 17776 44288
rect 17828 44276 17834 44328
rect 18509 44319 18567 44325
rect 18509 44285 18521 44319
rect 18555 44316 18567 44319
rect 19613 44319 19671 44325
rect 19613 44316 19625 44319
rect 18555 44288 19625 44316
rect 18555 44285 18567 44288
rect 18509 44279 18567 44285
rect 19613 44285 19625 44288
rect 19659 44285 19671 44319
rect 19613 44279 19671 44285
rect 19702 44276 19708 44328
rect 19760 44316 19766 44328
rect 19904 44316 19932 44356
rect 21910 44344 21916 44356
rect 21968 44344 21974 44396
rect 22002 44344 22008 44396
rect 22060 44384 22066 44396
rect 22097 44387 22155 44393
rect 22097 44384 22109 44387
rect 22060 44356 22109 44384
rect 22060 44344 22066 44356
rect 22097 44353 22109 44356
rect 22143 44353 22155 44387
rect 22204 44384 22232 44424
rect 22204 44356 22784 44384
rect 22097 44347 22155 44353
rect 19760 44288 19932 44316
rect 20533 44319 20591 44325
rect 19760 44276 19766 44288
rect 20533 44285 20545 44319
rect 20579 44316 20591 44319
rect 22554 44316 22560 44328
rect 20579 44288 22560 44316
rect 20579 44285 20591 44288
rect 20533 44279 20591 44285
rect 22554 44276 22560 44288
rect 22612 44276 22618 44328
rect 14001 44251 14059 44257
rect 12268 44220 13584 44248
rect 13648 44220 13860 44248
rect 11606 44140 11612 44192
rect 11664 44180 11670 44192
rect 13173 44183 13231 44189
rect 13173 44180 13185 44183
rect 11664 44152 13185 44180
rect 11664 44140 11670 44152
rect 13173 44149 13185 44152
rect 13219 44180 13231 44183
rect 13648 44180 13676 44220
rect 13219 44152 13676 44180
rect 13219 44149 13231 44152
rect 13173 44143 13231 44149
rect 13722 44140 13728 44192
rect 13780 44140 13786 44192
rect 13832 44180 13860 44220
rect 14001 44217 14013 44251
rect 14047 44248 14059 44251
rect 14090 44248 14096 44260
rect 14047 44220 14096 44248
rect 14047 44217 14059 44220
rect 14001 44211 14059 44217
rect 14090 44208 14096 44220
rect 14148 44208 14154 44260
rect 17586 44248 17592 44260
rect 14200 44220 14412 44248
rect 14200 44180 14228 44220
rect 13832 44152 14228 44180
rect 14384 44180 14412 44220
rect 15028 44220 17592 44248
rect 14734 44180 14740 44192
rect 14384 44152 14740 44180
rect 14734 44140 14740 44152
rect 14792 44140 14798 44192
rect 15028 44189 15056 44220
rect 17586 44208 17592 44220
rect 17644 44208 17650 44260
rect 17678 44208 17684 44260
rect 17736 44248 17742 44260
rect 18693 44251 18751 44257
rect 18693 44248 18705 44251
rect 17736 44220 18705 44248
rect 17736 44208 17742 44220
rect 18693 44217 18705 44220
rect 18739 44217 18751 44251
rect 18693 44211 18751 44217
rect 19061 44251 19119 44257
rect 19061 44217 19073 44251
rect 19107 44248 19119 44251
rect 20714 44248 20720 44260
rect 19107 44220 20720 44248
rect 19107 44217 19119 44220
rect 19061 44211 19119 44217
rect 20714 44208 20720 44220
rect 20772 44208 20778 44260
rect 21085 44251 21143 44257
rect 21085 44217 21097 44251
rect 21131 44248 21143 44251
rect 21913 44251 21971 44257
rect 21913 44248 21925 44251
rect 21131 44220 21925 44248
rect 21131 44217 21143 44220
rect 21085 44211 21143 44217
rect 21913 44217 21925 44220
rect 21959 44217 21971 44251
rect 21913 44211 21971 44217
rect 22649 44251 22707 44257
rect 22649 44217 22661 44251
rect 22695 44217 22707 44251
rect 22756 44248 22784 44356
rect 22940 44325 22968 44492
rect 26326 44480 26332 44492
rect 26384 44480 26390 44532
rect 26418 44480 26424 44532
rect 26476 44520 26482 44532
rect 26476 44492 32352 44520
rect 26476 44480 26482 44492
rect 23014 44412 23020 44464
rect 23072 44452 23078 44464
rect 27801 44455 27859 44461
rect 27801 44452 27813 44455
rect 23072 44424 27813 44452
rect 23072 44412 23078 44424
rect 27801 44421 27813 44424
rect 27847 44421 27859 44455
rect 31205 44455 31263 44461
rect 31205 44452 31217 44455
rect 27801 44415 27859 44421
rect 29840 44424 31217 44452
rect 23937 44387 23995 44393
rect 23937 44384 23949 44387
rect 23032 44356 23949 44384
rect 22925 44319 22983 44325
rect 22925 44285 22937 44319
rect 22971 44285 22983 44319
rect 22925 44279 22983 44285
rect 23032 44248 23060 44356
rect 23937 44353 23949 44356
rect 23983 44384 23995 44387
rect 24762 44384 24768 44396
rect 23983 44356 24768 44384
rect 23983 44353 23995 44356
rect 23937 44347 23995 44353
rect 24762 44344 24768 44356
rect 24820 44344 24826 44396
rect 24949 44387 25007 44393
rect 24949 44353 24961 44387
rect 24995 44384 25007 44387
rect 25038 44384 25044 44396
rect 24995 44356 25044 44384
rect 24995 44353 25007 44356
rect 24949 44347 25007 44353
rect 25038 44344 25044 44356
rect 25096 44344 25102 44396
rect 25682 44344 25688 44396
rect 25740 44344 25746 44396
rect 27338 44344 27344 44396
rect 27396 44384 27402 44396
rect 27617 44387 27675 44393
rect 27617 44384 27629 44387
rect 27396 44356 27629 44384
rect 27396 44344 27402 44356
rect 27617 44353 27629 44356
rect 27663 44353 27675 44387
rect 27617 44347 27675 44353
rect 28074 44344 28080 44396
rect 28132 44384 28138 44396
rect 28629 44387 28687 44393
rect 28629 44384 28641 44387
rect 28132 44356 28641 44384
rect 28132 44344 28138 44356
rect 28629 44353 28641 44356
rect 28675 44353 28687 44387
rect 28629 44347 28687 44353
rect 28718 44344 28724 44396
rect 28776 44384 28782 44396
rect 29840 44393 29868 44424
rect 31205 44421 31217 44424
rect 31251 44421 31263 44455
rect 32324 44452 32352 44492
rect 32398 44480 32404 44532
rect 32456 44480 32462 44532
rect 32950 44480 32956 44532
rect 33008 44520 33014 44532
rect 33008 44492 44496 44520
rect 33008 44480 33014 44492
rect 43438 44452 43444 44464
rect 32324 44424 38608 44452
rect 31205 44415 31263 44421
rect 28997 44387 29055 44393
rect 28997 44384 29009 44387
rect 28776 44356 29009 44384
rect 28776 44344 28782 44356
rect 28997 44353 29009 44356
rect 29043 44353 29055 44387
rect 28997 44347 29055 44353
rect 29825 44387 29883 44393
rect 29825 44353 29837 44387
rect 29871 44353 29883 44387
rect 29825 44347 29883 44353
rect 30377 44387 30435 44393
rect 30377 44353 30389 44387
rect 30423 44384 30435 44387
rect 30423 44356 32076 44384
rect 30423 44353 30435 44356
rect 30377 44347 30435 44353
rect 23109 44319 23167 44325
rect 23109 44285 23121 44319
rect 23155 44285 23167 44319
rect 23109 44279 23167 44285
rect 24121 44319 24179 44325
rect 24121 44285 24133 44319
rect 24167 44316 24179 44319
rect 27065 44319 27123 44325
rect 27065 44316 27077 44319
rect 24167 44288 27077 44316
rect 24167 44285 24179 44288
rect 24121 44279 24179 44285
rect 27065 44285 27077 44288
rect 27111 44285 27123 44319
rect 27065 44279 27123 44285
rect 22756 44220 23060 44248
rect 23124 44248 23152 44279
rect 27982 44276 27988 44328
rect 28040 44276 28046 44328
rect 31018 44276 31024 44328
rect 31076 44276 31082 44328
rect 32048 44325 32076 44356
rect 32600 44325 32628 44424
rect 33873 44387 33931 44393
rect 33873 44353 33885 44387
rect 33919 44384 33931 44387
rect 35158 44384 35164 44396
rect 33919 44356 35164 44384
rect 33919 44353 33931 44356
rect 33873 44347 33931 44353
rect 35158 44344 35164 44356
rect 35216 44344 35222 44396
rect 36909 44387 36967 44393
rect 36909 44353 36921 44387
rect 36955 44384 36967 44387
rect 38286 44384 38292 44396
rect 36955 44356 38292 44384
rect 36955 44353 36967 44356
rect 36909 44347 36967 44353
rect 38286 44344 38292 44356
rect 38344 44344 38350 44396
rect 31389 44319 31447 44325
rect 31389 44316 31401 44319
rect 31128 44288 31401 44316
rect 25222 44248 25228 44260
rect 23124 44220 25228 44248
rect 22649 44211 22707 44217
rect 15013 44183 15071 44189
rect 15013 44149 15025 44183
rect 15059 44149 15071 44183
rect 15013 44143 15071 44149
rect 15930 44140 15936 44192
rect 15988 44140 15994 44192
rect 16393 44183 16451 44189
rect 16393 44149 16405 44183
rect 16439 44180 16451 44183
rect 16850 44180 16856 44192
rect 16439 44152 16856 44180
rect 16439 44149 16451 44152
rect 16393 44143 16451 44149
rect 16850 44140 16856 44152
rect 16908 44140 16914 44192
rect 17773 44183 17831 44189
rect 17773 44149 17785 44183
rect 17819 44180 17831 44183
rect 18138 44180 18144 44192
rect 17819 44152 18144 44180
rect 17819 44149 17831 44152
rect 17773 44143 17831 44149
rect 18138 44140 18144 44152
rect 18196 44140 18202 44192
rect 18966 44140 18972 44192
rect 19024 44180 19030 44192
rect 19245 44183 19303 44189
rect 19245 44180 19257 44183
rect 19024 44152 19257 44180
rect 19024 44140 19030 44152
rect 19245 44149 19257 44152
rect 19291 44149 19303 44183
rect 19245 44143 19303 44149
rect 19705 44183 19763 44189
rect 19705 44149 19717 44183
rect 19751 44180 19763 44183
rect 19794 44180 19800 44192
rect 19751 44152 19800 44180
rect 19751 44149 19763 44152
rect 19705 44143 19763 44149
rect 19794 44140 19800 44152
rect 19852 44140 19858 44192
rect 21174 44140 21180 44192
rect 21232 44180 21238 44192
rect 21545 44183 21603 44189
rect 21545 44180 21557 44183
rect 21232 44152 21557 44180
rect 21232 44140 21238 44152
rect 21545 44149 21557 44152
rect 21591 44149 21603 44183
rect 21545 44143 21603 44149
rect 21726 44140 21732 44192
rect 21784 44180 21790 44192
rect 22005 44183 22063 44189
rect 22005 44180 22017 44183
rect 21784 44152 22017 44180
rect 21784 44140 21790 44152
rect 22005 44149 22017 44152
rect 22051 44149 22063 44183
rect 22664 44180 22692 44211
rect 25222 44208 25228 44220
rect 25280 44208 25286 44260
rect 25409 44251 25467 44257
rect 25409 44217 25421 44251
rect 25455 44248 25467 44251
rect 25498 44248 25504 44260
rect 25455 44220 25504 44248
rect 25455 44217 25467 44220
rect 25409 44211 25467 44217
rect 25498 44208 25504 44220
rect 25556 44208 25562 44260
rect 26878 44208 26884 44260
rect 26936 44208 26942 44260
rect 28445 44251 28503 44257
rect 28445 44217 28457 44251
rect 28491 44248 28503 44251
rect 30469 44251 30527 44257
rect 30469 44248 30481 44251
rect 28491 44220 30481 44248
rect 28491 44217 28503 44220
rect 28445 44211 28503 44217
rect 30469 44217 30481 44220
rect 30515 44217 30527 44251
rect 30469 44211 30527 44217
rect 23474 44180 23480 44192
rect 22664 44152 23480 44180
rect 22005 44143 22063 44149
rect 23474 44140 23480 44152
rect 23532 44140 23538 44192
rect 23658 44140 23664 44192
rect 23716 44140 23722 44192
rect 24210 44140 24216 44192
rect 24268 44180 24274 44192
rect 24305 44183 24363 44189
rect 24305 44180 24317 44183
rect 24268 44152 24317 44180
rect 24268 44140 24274 44152
rect 24305 44149 24317 44152
rect 24351 44149 24363 44183
rect 24305 44143 24363 44149
rect 24670 44140 24676 44192
rect 24728 44140 24734 44192
rect 24762 44140 24768 44192
rect 24820 44140 24826 44192
rect 25317 44183 25375 44189
rect 25317 44149 25329 44183
rect 25363 44180 25375 44183
rect 25682 44180 25688 44192
rect 25363 44152 25688 44180
rect 25363 44149 25375 44152
rect 25317 44143 25375 44149
rect 25682 44140 25688 44152
rect 25740 44140 25746 44192
rect 26237 44183 26295 44189
rect 26237 44149 26249 44183
rect 26283 44180 26295 44183
rect 26510 44180 26516 44192
rect 26283 44152 26516 44180
rect 26283 44149 26295 44152
rect 26237 44143 26295 44149
rect 26510 44140 26516 44152
rect 26568 44140 26574 44192
rect 27890 44140 27896 44192
rect 27948 44180 27954 44192
rect 28077 44183 28135 44189
rect 28077 44180 28089 44183
rect 27948 44152 28089 44180
rect 27948 44140 27954 44152
rect 28077 44149 28089 44152
rect 28123 44149 28135 44183
rect 28077 44143 28135 44149
rect 28537 44183 28595 44189
rect 28537 44149 28549 44183
rect 28583 44180 28595 44183
rect 28810 44180 28816 44192
rect 28583 44152 28816 44180
rect 28583 44149 28595 44152
rect 28537 44143 28595 44149
rect 28810 44140 28816 44152
rect 28868 44140 28874 44192
rect 29641 44183 29699 44189
rect 29641 44149 29653 44183
rect 29687 44180 29699 44183
rect 31128 44180 31156 44288
rect 31389 44285 31401 44288
rect 31435 44285 31447 44319
rect 31389 44279 31447 44285
rect 31849 44319 31907 44325
rect 31849 44285 31861 44319
rect 31895 44285 31907 44319
rect 31849 44279 31907 44285
rect 32033 44319 32091 44325
rect 32033 44285 32045 44319
rect 32079 44285 32091 44319
rect 32033 44279 32091 44285
rect 32217 44319 32275 44325
rect 32217 44285 32229 44319
rect 32263 44316 32275 44319
rect 32585 44319 32643 44325
rect 32585 44316 32597 44319
rect 32263 44288 32597 44316
rect 32263 44285 32275 44288
rect 32217 44279 32275 44285
rect 32585 44285 32597 44288
rect 32631 44285 32643 44319
rect 32585 44279 32643 44285
rect 31864 44248 31892 44279
rect 32232 44248 32260 44279
rect 33410 44276 33416 44328
rect 33468 44316 33474 44328
rect 34330 44316 34336 44328
rect 33468 44288 34336 44316
rect 33468 44276 33474 44288
rect 34330 44276 34336 44288
rect 34388 44316 34394 44328
rect 34701 44319 34759 44325
rect 34701 44316 34713 44319
rect 34388 44288 34713 44316
rect 34388 44276 34394 44288
rect 34701 44285 34713 44288
rect 34747 44285 34759 44319
rect 34701 44279 34759 44285
rect 35250 44276 35256 44328
rect 35308 44316 35314 44328
rect 35529 44319 35587 44325
rect 35529 44316 35541 44319
rect 35308 44288 35541 44316
rect 35308 44276 35314 44288
rect 35529 44285 35541 44288
rect 35575 44285 35587 44319
rect 35529 44279 35587 44285
rect 36722 44276 36728 44328
rect 36780 44316 36786 44328
rect 38580 44325 38608 44424
rect 40788 44424 43444 44452
rect 39393 44387 39451 44393
rect 39393 44353 39405 44387
rect 39439 44384 39451 44387
rect 39439 44356 39473 44384
rect 39439 44353 39451 44356
rect 39393 44347 39451 44353
rect 38105 44319 38163 44325
rect 38105 44316 38117 44319
rect 36780 44288 38117 44316
rect 36780 44276 36786 44288
rect 38105 44285 38117 44288
rect 38151 44285 38163 44319
rect 38105 44279 38163 44285
rect 38565 44319 38623 44325
rect 38565 44285 38577 44319
rect 38611 44285 38623 44319
rect 38565 44279 38623 44285
rect 38838 44276 38844 44328
rect 38896 44276 38902 44328
rect 39408 44316 39436 44347
rect 39942 44316 39948 44328
rect 39224 44288 39948 44316
rect 33318 44248 33324 44260
rect 31864 44220 32260 44248
rect 33152 44220 33324 44248
rect 29687 44152 31156 44180
rect 29687 44149 29699 44152
rect 29641 44143 29699 44149
rect 31294 44140 31300 44192
rect 31352 44180 31358 44192
rect 31665 44183 31723 44189
rect 31665 44180 31677 44183
rect 31352 44152 31677 44180
rect 31352 44140 31358 44152
rect 31665 44149 31677 44152
rect 31711 44180 31723 44183
rect 33152 44180 33180 44220
rect 33318 44208 33324 44220
rect 33376 44208 33382 44260
rect 33597 44251 33655 44257
rect 33597 44217 33609 44251
rect 33643 44248 33655 44251
rect 34149 44251 34207 44257
rect 34149 44248 34161 44251
rect 33643 44220 34161 44248
rect 33643 44217 33655 44220
rect 33597 44211 33655 44217
rect 34149 44217 34161 44220
rect 34195 44217 34207 44251
rect 36081 44251 36139 44257
rect 36081 44248 36093 44251
rect 34149 44211 34207 44217
rect 35544 44220 36093 44248
rect 35544 44192 35572 44220
rect 36081 44217 36093 44220
rect 36127 44217 36139 44251
rect 36081 44211 36139 44217
rect 37093 44251 37151 44257
rect 37093 44217 37105 44251
rect 37139 44248 37151 44251
rect 37553 44251 37611 44257
rect 37553 44248 37565 44251
rect 37139 44220 37565 44248
rect 37139 44217 37151 44220
rect 37093 44211 37151 44217
rect 37553 44217 37565 44220
rect 37599 44217 37611 44251
rect 37553 44211 37611 44217
rect 37734 44208 37740 44260
rect 37792 44248 37798 44260
rect 39224 44248 39252 44288
rect 39942 44276 39948 44288
rect 40000 44276 40006 44328
rect 40310 44276 40316 44328
rect 40368 44316 40374 44328
rect 40497 44319 40555 44325
rect 40497 44316 40509 44319
rect 40368 44288 40509 44316
rect 40368 44276 40374 44288
rect 40497 44285 40509 44288
rect 40543 44285 40555 44319
rect 40497 44279 40555 44285
rect 37792 44220 39252 44248
rect 37792 44208 37798 44220
rect 39298 44208 39304 44260
rect 39356 44248 39362 44260
rect 39669 44251 39727 44257
rect 39669 44248 39681 44251
rect 39356 44220 39681 44248
rect 39356 44208 39362 44220
rect 39669 44217 39681 44220
rect 39715 44248 39727 44251
rect 40788 44248 40816 44424
rect 43438 44412 43444 44424
rect 43496 44412 43502 44464
rect 41414 44344 41420 44396
rect 41472 44384 41478 44396
rect 42429 44387 42487 44393
rect 42429 44384 42441 44387
rect 41472 44356 42441 44384
rect 41472 44344 41478 44356
rect 42429 44353 42441 44356
rect 42475 44353 42487 44387
rect 44358 44384 44364 44396
rect 42429 44347 42487 44353
rect 42904 44356 44364 44384
rect 41049 44319 41107 44325
rect 41049 44285 41061 44319
rect 41095 44316 41107 44319
rect 41230 44316 41236 44328
rect 41095 44288 41236 44316
rect 41095 44285 41107 44288
rect 41049 44279 41107 44285
rect 41230 44276 41236 44288
rect 41288 44316 41294 44328
rect 42904 44316 42932 44356
rect 44358 44344 44364 44356
rect 44416 44344 44422 44396
rect 41288 44288 42932 44316
rect 41288 44276 41294 44288
rect 43346 44276 43352 44328
rect 43404 44276 43410 44328
rect 44085 44319 44143 44325
rect 44085 44285 44097 44319
rect 44131 44316 44143 44319
rect 44174 44316 44180 44328
rect 44131 44288 44180 44316
rect 44131 44285 44143 44288
rect 44085 44279 44143 44285
rect 44174 44276 44180 44288
rect 44232 44276 44238 44328
rect 44468 44325 44496 44492
rect 46661 44455 46719 44461
rect 46661 44421 46673 44455
rect 46707 44452 46719 44455
rect 47394 44452 47400 44464
rect 46707 44424 47400 44452
rect 46707 44421 46719 44424
rect 46661 44415 46719 44421
rect 47394 44412 47400 44424
rect 47452 44412 47458 44464
rect 46106 44344 46112 44396
rect 46164 44384 46170 44396
rect 46293 44387 46351 44393
rect 46293 44384 46305 44387
rect 46164 44356 46305 44384
rect 46164 44344 46170 44356
rect 46293 44353 46305 44356
rect 46339 44353 46351 44387
rect 46293 44347 46351 44353
rect 44453 44319 44511 44325
rect 44453 44285 44465 44319
rect 44499 44285 44511 44319
rect 44453 44279 44511 44285
rect 45922 44276 45928 44328
rect 45980 44316 45986 44328
rect 46201 44319 46259 44325
rect 46201 44316 46213 44319
rect 45980 44288 46213 44316
rect 45980 44276 45986 44288
rect 46201 44285 46213 44288
rect 46247 44285 46259 44319
rect 46201 44279 46259 44285
rect 46845 44319 46903 44325
rect 46845 44285 46857 44319
rect 46891 44316 46903 44319
rect 52730 44316 52736 44328
rect 46891 44288 52736 44316
rect 46891 44285 46903 44288
rect 46845 44279 46903 44285
rect 52730 44276 52736 44288
rect 52788 44276 52794 44328
rect 41325 44251 41383 44257
rect 41325 44248 41337 44251
rect 39715 44220 40816 44248
rect 40972 44220 41337 44248
rect 39715 44217 39727 44220
rect 39669 44211 39727 44217
rect 31711 44152 33180 44180
rect 31711 44149 31723 44152
rect 31665 44143 31723 44149
rect 33226 44140 33232 44192
rect 33284 44140 33290 44192
rect 33689 44183 33747 44189
rect 33689 44149 33701 44183
rect 33735 44180 33747 44183
rect 34422 44180 34428 44192
rect 33735 44152 34428 44180
rect 33735 44149 33747 44152
rect 33689 44143 33747 44149
rect 34422 44140 34428 44152
rect 34480 44140 34486 44192
rect 34514 44140 34520 44192
rect 34572 44180 34578 44192
rect 34977 44183 35035 44189
rect 34977 44180 34989 44183
rect 34572 44152 34989 44180
rect 34572 44140 34578 44152
rect 34977 44149 34989 44152
rect 35023 44149 35035 44183
rect 34977 44143 35035 44149
rect 35526 44140 35532 44192
rect 35584 44140 35590 44192
rect 35802 44140 35808 44192
rect 35860 44140 35866 44192
rect 36538 44140 36544 44192
rect 36596 44180 36602 44192
rect 37001 44183 37059 44189
rect 37001 44180 37013 44183
rect 36596 44152 37013 44180
rect 36596 44140 36602 44152
rect 37001 44149 37013 44152
rect 37047 44149 37059 44183
rect 37001 44143 37059 44149
rect 37461 44183 37519 44189
rect 37461 44149 37473 44183
rect 37507 44180 37519 44183
rect 38194 44180 38200 44192
rect 37507 44152 38200 44180
rect 37507 44149 37519 44152
rect 37461 44143 37519 44149
rect 38194 44140 38200 44152
rect 38252 44140 38258 44192
rect 39482 44140 39488 44192
rect 39540 44180 39546 44192
rect 39945 44183 40003 44189
rect 39945 44180 39957 44183
rect 39540 44152 39957 44180
rect 39540 44140 39546 44152
rect 39945 44149 39957 44152
rect 39991 44149 40003 44183
rect 39945 44143 40003 44149
rect 40862 44140 40868 44192
rect 40920 44180 40926 44192
rect 40972 44189 41000 44220
rect 41325 44217 41337 44220
rect 41371 44217 41383 44251
rect 41325 44211 41383 44217
rect 42245 44251 42303 44257
rect 42245 44217 42257 44251
rect 42291 44248 42303 44251
rect 43441 44251 43499 44257
rect 43441 44248 43453 44251
rect 42291 44220 43453 44248
rect 42291 44217 42303 44220
rect 42245 44211 42303 44217
rect 43441 44217 43453 44220
rect 43487 44217 43499 44251
rect 43441 44211 43499 44217
rect 44726 44208 44732 44260
rect 44784 44248 44790 44260
rect 44784 44220 47256 44248
rect 44784 44208 44790 44220
rect 40957 44183 41015 44189
rect 40957 44180 40969 44183
rect 40920 44152 40969 44180
rect 40920 44140 40926 44152
rect 40957 44149 40969 44152
rect 41003 44149 41015 44183
rect 40957 44143 41015 44149
rect 41414 44140 41420 44192
rect 41472 44140 41478 44192
rect 41877 44183 41935 44189
rect 41877 44149 41889 44183
rect 41923 44180 41935 44183
rect 42150 44180 42156 44192
rect 41923 44152 42156 44180
rect 41923 44149 41935 44152
rect 41877 44143 41935 44149
rect 42150 44140 42156 44152
rect 42208 44140 42214 44192
rect 42334 44140 42340 44192
rect 42392 44140 42398 44192
rect 42518 44140 42524 44192
rect 42576 44180 42582 44192
rect 42705 44183 42763 44189
rect 42705 44180 42717 44183
rect 42576 44152 42717 44180
rect 42576 44140 42582 44152
rect 42705 44149 42717 44152
rect 42751 44149 42763 44183
rect 42705 44143 42763 44149
rect 45370 44140 45376 44192
rect 45428 44180 45434 44192
rect 45741 44183 45799 44189
rect 45741 44180 45753 44183
rect 45428 44152 45753 44180
rect 45428 44140 45434 44152
rect 45741 44149 45753 44152
rect 45787 44149 45799 44183
rect 45741 44143 45799 44149
rect 46014 44140 46020 44192
rect 46072 44180 46078 44192
rect 46109 44183 46167 44189
rect 46109 44180 46121 44183
rect 46072 44152 46121 44180
rect 46072 44140 46078 44152
rect 46109 44149 46121 44152
rect 46155 44149 46167 44183
rect 46109 44143 46167 44149
rect 46658 44140 46664 44192
rect 46716 44180 46722 44192
rect 47121 44183 47179 44189
rect 47121 44180 47133 44183
rect 46716 44152 47133 44180
rect 46716 44140 46722 44152
rect 47121 44149 47133 44152
rect 47167 44149 47179 44183
rect 47228 44180 47256 44220
rect 47394 44208 47400 44260
rect 47452 44248 47458 44260
rect 48038 44248 48044 44260
rect 47452 44220 48044 44248
rect 47452 44208 47458 44220
rect 48038 44208 48044 44220
rect 48096 44208 48102 44260
rect 53834 44180 53840 44192
rect 47228 44152 53840 44180
rect 47121 44143 47179 44149
rect 53834 44140 53840 44152
rect 53892 44140 53898 44192
rect 552 44090 66424 44112
rect 552 44038 2918 44090
rect 2970 44038 2982 44090
rect 3034 44038 3046 44090
rect 3098 44038 3110 44090
rect 3162 44038 3174 44090
rect 3226 44038 50918 44090
rect 50970 44038 50982 44090
rect 51034 44038 51046 44090
rect 51098 44038 51110 44090
rect 51162 44038 51174 44090
rect 51226 44038 66424 44090
rect 552 44016 66424 44038
rect 14001 43979 14059 43985
rect 14001 43945 14013 43979
rect 14047 43976 14059 43979
rect 14642 43976 14648 43988
rect 14047 43948 14648 43976
rect 14047 43945 14059 43948
rect 14001 43939 14059 43945
rect 14642 43936 14648 43948
rect 14700 43976 14706 43988
rect 14700 43948 15884 43976
rect 14700 43936 14706 43948
rect 11517 43911 11575 43917
rect 11517 43877 11529 43911
rect 11563 43908 11575 43911
rect 12526 43908 12532 43920
rect 11563 43880 12532 43908
rect 11563 43877 11575 43880
rect 11517 43871 11575 43877
rect 12526 43868 12532 43880
rect 12584 43868 12590 43920
rect 12897 43911 12955 43917
rect 12897 43877 12909 43911
rect 12943 43908 12955 43911
rect 13449 43911 13507 43917
rect 13449 43908 13461 43911
rect 12943 43880 13461 43908
rect 12943 43877 12955 43880
rect 12897 43871 12955 43877
rect 13449 43877 13461 43880
rect 13495 43877 13507 43911
rect 13449 43871 13507 43877
rect 11425 43843 11483 43849
rect 11425 43809 11437 43843
rect 11471 43840 11483 43843
rect 11885 43843 11943 43849
rect 11885 43840 11897 43843
rect 11471 43812 11897 43840
rect 11471 43809 11483 43812
rect 11425 43803 11483 43809
rect 11885 43809 11897 43812
rect 11931 43809 11943 43843
rect 11885 43803 11943 43809
rect 12802 43800 12808 43852
rect 12860 43800 12866 43852
rect 11606 43732 11612 43784
rect 11664 43732 11670 43784
rect 11698 43732 11704 43784
rect 11756 43772 11762 43784
rect 12437 43775 12495 43781
rect 12437 43772 12449 43775
rect 11756 43744 12449 43772
rect 11756 43732 11762 43744
rect 12437 43741 12449 43744
rect 12483 43741 12495 43775
rect 12437 43735 12495 43741
rect 12250 43664 12256 43716
rect 12308 43704 12314 43716
rect 12912 43704 12940 43871
rect 13722 43868 13728 43920
rect 13780 43908 13786 43920
rect 14093 43911 14151 43917
rect 14093 43908 14105 43911
rect 13780 43880 14105 43908
rect 13780 43868 13786 43880
rect 14093 43877 14105 43880
rect 14139 43877 14151 43911
rect 14093 43871 14151 43877
rect 14921 43911 14979 43917
rect 14921 43877 14933 43911
rect 14967 43908 14979 43911
rect 15194 43908 15200 43920
rect 14967 43880 15200 43908
rect 14967 43877 14979 43880
rect 14921 43871 14979 43877
rect 15194 43868 15200 43880
rect 15252 43868 15258 43920
rect 15856 43849 15884 43948
rect 15930 43936 15936 43988
rect 15988 43976 15994 43988
rect 16853 43979 16911 43985
rect 16853 43976 16865 43979
rect 15988 43948 16865 43976
rect 15988 43936 15994 43948
rect 16853 43945 16865 43948
rect 16899 43945 16911 43979
rect 16853 43939 16911 43945
rect 16945 43979 17003 43985
rect 16945 43945 16957 43979
rect 16991 43976 17003 43979
rect 17313 43979 17371 43985
rect 17313 43976 17325 43979
rect 16991 43948 17325 43976
rect 16991 43945 17003 43948
rect 16945 43939 17003 43945
rect 17313 43945 17325 43948
rect 17359 43945 17371 43979
rect 17313 43939 17371 43945
rect 17402 43936 17408 43988
rect 17460 43976 17466 43988
rect 17681 43979 17739 43985
rect 17681 43976 17693 43979
rect 17460 43948 17693 43976
rect 17460 43936 17466 43948
rect 17681 43945 17693 43948
rect 17727 43945 17739 43979
rect 17681 43939 17739 43945
rect 17770 43936 17776 43988
rect 17828 43936 17834 43988
rect 18322 43936 18328 43988
rect 18380 43936 18386 43988
rect 20714 43976 20720 43988
rect 20456 43948 20720 43976
rect 17788 43908 17816 43936
rect 19334 43908 19340 43920
rect 17052 43880 17540 43908
rect 17788 43880 19340 43908
rect 13081 43843 13139 43849
rect 13081 43809 13093 43843
rect 13127 43840 13139 43843
rect 14829 43843 14887 43849
rect 13127 43812 14780 43840
rect 13127 43809 13139 43812
rect 13081 43803 13139 43809
rect 14185 43775 14243 43781
rect 12308 43676 12940 43704
rect 13004 43744 13952 43772
rect 12308 43664 12314 43676
rect 11054 43596 11060 43648
rect 11112 43596 11118 43648
rect 12618 43596 12624 43648
rect 12676 43636 12682 43648
rect 13004 43636 13032 43744
rect 13265 43707 13323 43713
rect 13265 43673 13277 43707
rect 13311 43704 13323 43707
rect 13814 43704 13820 43716
rect 13311 43676 13820 43704
rect 13311 43673 13323 43676
rect 13265 43667 13323 43673
rect 13814 43664 13820 43676
rect 13872 43664 13878 43716
rect 13924 43704 13952 43744
rect 14185 43741 14197 43775
rect 14231 43741 14243 43775
rect 14185 43735 14243 43741
rect 14200 43704 14228 43735
rect 13924 43676 14228 43704
rect 14752 43704 14780 43812
rect 14829 43809 14841 43843
rect 14875 43840 14887 43843
rect 15289 43843 15347 43849
rect 15289 43840 15301 43843
rect 14875 43812 15301 43840
rect 14875 43809 14887 43812
rect 14829 43803 14887 43809
rect 15289 43809 15301 43812
rect 15335 43809 15347 43843
rect 15289 43803 15347 43809
rect 15841 43843 15899 43849
rect 15841 43809 15853 43843
rect 15887 43809 15899 43843
rect 15841 43803 15899 43809
rect 16206 43800 16212 43852
rect 16264 43800 16270 43852
rect 14918 43732 14924 43784
rect 14976 43772 14982 43784
rect 15013 43775 15071 43781
rect 15013 43772 15025 43775
rect 14976 43744 15025 43772
rect 14976 43732 14982 43744
rect 15013 43741 15025 43744
rect 15059 43741 15071 43775
rect 15013 43735 15071 43741
rect 17052 43704 17080 43880
rect 17129 43775 17187 43781
rect 17129 43741 17141 43775
rect 17175 43772 17187 43775
rect 17175 43744 17356 43772
rect 17175 43741 17187 43744
rect 17129 43735 17187 43741
rect 14752 43676 17080 43704
rect 12676 43608 13032 43636
rect 12676 43596 12682 43608
rect 13630 43596 13636 43648
rect 13688 43596 13694 43648
rect 14458 43596 14464 43648
rect 14516 43596 14522 43648
rect 15930 43596 15936 43648
rect 15988 43636 15994 43648
rect 16485 43639 16543 43645
rect 16485 43636 16497 43639
rect 15988 43608 16497 43636
rect 15988 43596 15994 43608
rect 16485 43605 16497 43608
rect 16531 43605 16543 43639
rect 16485 43599 16543 43605
rect 17126 43596 17132 43648
rect 17184 43636 17190 43648
rect 17328 43636 17356 43744
rect 17512 43704 17540 43880
rect 19334 43868 19340 43880
rect 19392 43868 19398 43920
rect 20456 43908 20484 43948
rect 20714 43936 20720 43948
rect 20772 43976 20778 43988
rect 21542 43976 21548 43988
rect 20772 43948 21548 43976
rect 20772 43936 20778 43948
rect 21542 43936 21548 43948
rect 21600 43936 21606 43988
rect 21726 43936 21732 43988
rect 21784 43936 21790 43988
rect 23937 43979 23995 43985
rect 23937 43945 23949 43979
rect 23983 43976 23995 43979
rect 24670 43976 24676 43988
rect 23983 43948 24676 43976
rect 23983 43945 23995 43948
rect 23937 43939 23995 43945
rect 24670 43936 24676 43948
rect 24728 43936 24734 43988
rect 24946 43936 24952 43988
rect 25004 43976 25010 43988
rect 32950 43976 32956 43988
rect 25004 43948 32956 43976
rect 25004 43936 25010 43948
rect 20378 43880 20484 43908
rect 20809 43911 20867 43917
rect 20809 43877 20821 43911
rect 20855 43908 20867 43911
rect 20855 43880 21864 43908
rect 20855 43877 20867 43880
rect 20809 43871 20867 43877
rect 18509 43843 18567 43849
rect 18509 43809 18521 43843
rect 18555 43840 18567 43843
rect 18693 43843 18751 43849
rect 18693 43840 18705 43843
rect 18555 43812 18705 43840
rect 18555 43809 18567 43812
rect 18509 43803 18567 43809
rect 18693 43809 18705 43812
rect 18739 43840 18751 43843
rect 19426 43840 19432 43852
rect 18739 43812 19432 43840
rect 18739 43809 18751 43812
rect 18693 43803 18751 43809
rect 19426 43800 19432 43812
rect 19484 43800 19490 43852
rect 21634 43800 21640 43852
rect 21692 43800 21698 43852
rect 21836 43840 21864 43880
rect 21910 43868 21916 43920
rect 21968 43908 21974 43920
rect 22097 43911 22155 43917
rect 22097 43908 22109 43911
rect 21968 43880 22109 43908
rect 21968 43868 21974 43880
rect 22097 43877 22109 43880
rect 22143 43877 22155 43911
rect 22097 43871 22155 43877
rect 22189 43911 22247 43917
rect 22189 43877 22201 43911
rect 22235 43908 22247 43911
rect 23014 43908 23020 43920
rect 22235 43880 23020 43908
rect 22235 43877 22247 43880
rect 22189 43871 22247 43877
rect 23014 43868 23020 43880
rect 23072 43868 23078 43920
rect 23658 43868 23664 43920
rect 23716 43908 23722 43920
rect 24305 43911 24363 43917
rect 24305 43908 24317 43911
rect 23716 43880 24317 43908
rect 23716 43868 23722 43880
rect 24305 43877 24317 43880
rect 24351 43877 24363 43911
rect 24305 43871 24363 43877
rect 24854 43868 24860 43920
rect 24912 43868 24918 43920
rect 26160 43917 26188 43948
rect 32950 43936 32956 43948
rect 33008 43936 33014 43988
rect 33410 43936 33416 43988
rect 33468 43936 33474 43988
rect 36538 43936 36544 43988
rect 36596 43936 36602 43988
rect 36722 43936 36728 43988
rect 36780 43936 36786 43988
rect 36924 43948 39160 43976
rect 26145 43911 26203 43917
rect 26145 43877 26157 43911
rect 26191 43877 26203 43911
rect 26145 43871 26203 43877
rect 27617 43911 27675 43917
rect 27617 43877 27629 43911
rect 27663 43908 27675 43911
rect 27890 43908 27896 43920
rect 27663 43880 27896 43908
rect 27663 43877 27675 43880
rect 27617 43871 27675 43877
rect 27890 43868 27896 43880
rect 27948 43868 27954 43920
rect 29086 43908 29092 43920
rect 28842 43880 29092 43908
rect 29086 43868 29092 43880
rect 29144 43868 29150 43920
rect 32214 43908 32220 43920
rect 31680 43880 32220 43908
rect 22278 43840 22284 43852
rect 21836 43812 22284 43840
rect 22278 43800 22284 43812
rect 22336 43800 22342 43852
rect 26234 43800 26240 43852
rect 26292 43840 26298 43852
rect 26878 43840 26884 43852
rect 26292 43812 26884 43840
rect 26292 43800 26298 43812
rect 26878 43800 26884 43812
rect 26936 43840 26942 43852
rect 27341 43843 27399 43849
rect 27341 43840 27353 43843
rect 26936 43812 27353 43840
rect 26936 43800 26942 43812
rect 27341 43809 27353 43812
rect 27387 43809 27399 43843
rect 27341 43803 27399 43809
rect 30558 43800 30564 43852
rect 30616 43800 30622 43852
rect 31680 43849 31708 43880
rect 32214 43868 32220 43880
rect 32272 43868 32278 43920
rect 33318 43908 33324 43920
rect 33166 43880 33324 43908
rect 33318 43868 33324 43880
rect 33376 43908 33382 43920
rect 33376 43880 34270 43908
rect 33376 43868 33382 43880
rect 35250 43868 35256 43920
rect 35308 43908 35314 43920
rect 36081 43911 36139 43917
rect 36081 43908 36093 43911
rect 35308 43880 36093 43908
rect 35308 43868 35314 43880
rect 36081 43877 36093 43880
rect 36127 43877 36139 43911
rect 36081 43871 36139 43877
rect 36173 43911 36231 43917
rect 36173 43877 36185 43911
rect 36219 43908 36231 43911
rect 36354 43908 36360 43920
rect 36219 43880 36360 43908
rect 36219 43877 36231 43880
rect 36173 43871 36231 43877
rect 36354 43868 36360 43880
rect 36412 43908 36418 43920
rect 36924 43908 36952 43948
rect 36412 43880 36952 43908
rect 36412 43868 36418 43880
rect 37734 43868 37740 43920
rect 37792 43868 37798 43920
rect 38194 43868 38200 43920
rect 38252 43868 38258 43920
rect 31665 43843 31723 43849
rect 31665 43809 31677 43843
rect 31711 43809 31723 43843
rect 31665 43803 31723 43809
rect 35434 43800 35440 43852
rect 35492 43800 35498 43852
rect 39132 43849 39160 43948
rect 39390 43936 39396 43988
rect 39448 43976 39454 43988
rect 39485 43979 39543 43985
rect 39485 43976 39497 43979
rect 39448 43948 39497 43976
rect 39448 43936 39454 43948
rect 39485 43945 39497 43948
rect 39531 43945 39543 43979
rect 39485 43939 39543 43945
rect 41230 43936 41236 43988
rect 41288 43976 41294 43988
rect 41417 43979 41475 43985
rect 41417 43976 41429 43979
rect 41288 43948 41429 43976
rect 41288 43936 41294 43948
rect 41417 43945 41429 43948
rect 41463 43945 41475 43979
rect 44726 43976 44732 43988
rect 41417 43939 41475 43945
rect 41524 43948 44732 43976
rect 41524 43917 41552 43948
rect 44726 43936 44732 43948
rect 44784 43936 44790 43988
rect 46845 43979 46903 43985
rect 46845 43945 46857 43979
rect 46891 43976 46903 43979
rect 47397 43979 47455 43985
rect 47397 43976 47409 43979
rect 46891 43948 47409 43976
rect 46891 43945 46903 43948
rect 46845 43939 46903 43945
rect 47397 43945 47409 43948
rect 47443 43945 47455 43979
rect 47397 43939 47455 43945
rect 41509 43911 41567 43917
rect 40526 43880 41414 43908
rect 39117 43843 39175 43849
rect 39117 43809 39129 43843
rect 39163 43809 39175 43843
rect 39117 43803 39175 43809
rect 17586 43732 17592 43784
rect 17644 43772 17650 43784
rect 17862 43772 17868 43784
rect 17644 43744 17868 43772
rect 17644 43732 17650 43744
rect 17862 43732 17868 43744
rect 17920 43732 17926 43784
rect 19245 43775 19303 43781
rect 19245 43741 19257 43775
rect 19291 43772 19303 43775
rect 19291 43744 21036 43772
rect 19291 43741 19303 43744
rect 19245 43735 19303 43741
rect 21008 43704 21036 43744
rect 21082 43732 21088 43784
rect 21140 43732 21146 43784
rect 22094 43772 22100 43784
rect 21192 43744 22100 43772
rect 21192 43704 21220 43744
rect 22094 43732 22100 43744
rect 22152 43732 22158 43784
rect 22370 43732 22376 43784
rect 22428 43732 22434 43784
rect 22738 43732 22744 43784
rect 22796 43772 22802 43784
rect 23109 43775 23167 43781
rect 23109 43772 23121 43775
rect 22796 43744 23121 43772
rect 22796 43732 22802 43744
rect 23109 43741 23121 43744
rect 23155 43741 23167 43775
rect 23109 43735 23167 43741
rect 23382 43732 23388 43784
rect 23440 43732 23446 43784
rect 24029 43775 24087 43781
rect 24029 43741 24041 43775
rect 24075 43772 24087 43775
rect 26421 43775 26479 43781
rect 24075 43744 26372 43772
rect 24075 43741 24087 43744
rect 24029 43735 24087 43741
rect 17512 43676 19840 43704
rect 21008 43676 21220 43704
rect 18414 43636 18420 43648
rect 17184 43608 18420 43636
rect 17184 43596 17190 43608
rect 18414 43596 18420 43608
rect 18472 43596 18478 43648
rect 19337 43639 19395 43645
rect 19337 43605 19349 43639
rect 19383 43636 19395 43639
rect 19426 43636 19432 43648
rect 19383 43608 19432 43636
rect 19383 43605 19395 43608
rect 19337 43599 19395 43605
rect 19426 43596 19432 43608
rect 19484 43636 19490 43648
rect 19702 43636 19708 43648
rect 19484 43608 19708 43636
rect 19484 43596 19490 43608
rect 19702 43596 19708 43608
rect 19760 43596 19766 43648
rect 19812 43636 19840 43676
rect 21450 43664 21456 43716
rect 21508 43704 21514 43716
rect 21818 43704 21824 43716
rect 21508 43676 21824 43704
rect 21508 43664 21514 43676
rect 21818 43664 21824 43676
rect 21876 43664 21882 43716
rect 26344 43704 26372 43744
rect 26421 43741 26433 43775
rect 26467 43772 26479 43775
rect 26786 43772 26792 43784
rect 26467 43744 26792 43772
rect 26467 43741 26479 43744
rect 26421 43735 26479 43741
rect 26786 43732 26792 43744
rect 26844 43732 26850 43784
rect 27065 43775 27123 43781
rect 27065 43741 27077 43775
rect 27111 43772 27123 43775
rect 27246 43772 27252 43784
rect 27111 43744 27252 43772
rect 27111 43741 27123 43744
rect 27065 43735 27123 43741
rect 27246 43732 27252 43744
rect 27304 43732 27310 43784
rect 29181 43775 29239 43781
rect 29181 43772 29193 43775
rect 27356 43744 29193 43772
rect 26602 43704 26608 43716
rect 26344 43676 26608 43704
rect 26602 43664 26608 43676
rect 26660 43704 26666 43716
rect 27356 43704 27384 43744
rect 29181 43741 29193 43744
rect 29227 43741 29239 43775
rect 29181 43735 29239 43741
rect 29457 43775 29515 43781
rect 29457 43741 29469 43775
rect 29503 43772 29515 43775
rect 29546 43772 29552 43784
rect 29503 43744 29552 43772
rect 29503 43741 29515 43744
rect 29457 43735 29515 43741
rect 29546 43732 29552 43744
rect 29604 43732 29610 43784
rect 29914 43732 29920 43784
rect 29972 43772 29978 43784
rect 31205 43775 31263 43781
rect 31205 43772 31217 43775
rect 29972 43744 31217 43772
rect 29972 43732 29978 43744
rect 31205 43741 31217 43744
rect 31251 43741 31263 43775
rect 31205 43735 31263 43741
rect 31941 43775 31999 43781
rect 31941 43741 31953 43775
rect 31987 43772 31999 43775
rect 33226 43772 33232 43784
rect 31987 43744 33232 43772
rect 31987 43741 31999 43744
rect 31941 43735 31999 43741
rect 33226 43732 33232 43744
rect 33284 43732 33290 43784
rect 33505 43775 33563 43781
rect 33505 43741 33517 43775
rect 33551 43772 33563 43775
rect 33781 43775 33839 43781
rect 33551 43744 33640 43772
rect 33551 43741 33563 43744
rect 33505 43735 33563 43741
rect 26660 43676 27384 43704
rect 26660 43664 26666 43676
rect 20070 43636 20076 43648
rect 19812 43608 20076 43636
rect 20070 43596 20076 43608
rect 20128 43596 20134 43648
rect 20162 43596 20168 43648
rect 20220 43636 20226 43648
rect 21082 43636 21088 43648
rect 20220 43608 21088 43636
rect 20220 43596 20226 43608
rect 21082 43596 21088 43608
rect 21140 43596 21146 43648
rect 22462 43596 22468 43648
rect 22520 43636 22526 43648
rect 22557 43639 22615 43645
rect 22557 43636 22569 43639
rect 22520 43608 22569 43636
rect 22520 43596 22526 43608
rect 22557 43605 22569 43608
rect 22603 43605 22615 43639
rect 22557 43599 22615 43605
rect 25777 43639 25835 43645
rect 25777 43605 25789 43639
rect 25823 43636 25835 43639
rect 25866 43636 25872 43648
rect 25823 43608 25872 43636
rect 25823 43605 25835 43608
rect 25777 43599 25835 43605
rect 25866 43596 25872 43608
rect 25924 43596 25930 43648
rect 26050 43596 26056 43648
rect 26108 43596 26114 43648
rect 29089 43639 29147 43645
rect 29089 43605 29101 43639
rect 29135 43636 29147 43639
rect 31018 43636 31024 43648
rect 29135 43608 31024 43636
rect 29135 43605 29147 43608
rect 29089 43599 29147 43605
rect 31018 43596 31024 43608
rect 31076 43596 31082 43648
rect 31754 43596 31760 43648
rect 31812 43636 31818 43648
rect 33612 43636 33640 43744
rect 33781 43741 33793 43775
rect 33827 43772 33839 43775
rect 34146 43772 34152 43784
rect 33827 43744 34152 43772
rect 33827 43741 33839 43744
rect 33781 43735 33839 43741
rect 34146 43732 34152 43744
rect 34204 43732 34210 43784
rect 35342 43732 35348 43784
rect 35400 43772 35406 43784
rect 35802 43772 35808 43784
rect 35400 43744 35808 43772
rect 35400 43732 35406 43744
rect 35802 43732 35808 43744
rect 35860 43772 35866 43784
rect 35897 43775 35955 43781
rect 35897 43772 35909 43775
rect 35860 43744 35909 43772
rect 35860 43732 35866 43744
rect 35897 43741 35909 43744
rect 35943 43741 35955 43775
rect 35897 43735 35955 43741
rect 38470 43732 38476 43784
rect 38528 43732 38534 43784
rect 40954 43732 40960 43784
rect 41012 43732 41018 43784
rect 41230 43732 41236 43784
rect 41288 43732 41294 43784
rect 41386 43704 41414 43880
rect 41509 43877 41521 43911
rect 41555 43877 41567 43911
rect 41509 43871 41567 43877
rect 42150 43868 42156 43920
rect 42208 43868 42214 43920
rect 43438 43868 43444 43920
rect 43496 43908 43502 43920
rect 44453 43911 44511 43917
rect 44453 43908 44465 43911
rect 43496 43880 44465 43908
rect 43496 43868 43502 43880
rect 44453 43877 44465 43880
rect 44499 43877 44511 43911
rect 46658 43908 46664 43920
rect 46598 43880 46664 43908
rect 44453 43871 44511 43877
rect 46658 43868 46664 43880
rect 46716 43868 46722 43920
rect 41874 43732 41880 43784
rect 41932 43732 41938 43784
rect 43162 43772 43168 43784
rect 41984 43744 43168 43772
rect 41984 43704 42012 43744
rect 43162 43732 43168 43744
rect 43220 43772 43226 43784
rect 43272 43772 43300 43826
rect 43898 43800 43904 43852
rect 43956 43840 43962 43852
rect 44085 43843 44143 43849
rect 44085 43840 44097 43843
rect 43956 43812 44097 43840
rect 43956 43800 43962 43812
rect 44085 43809 44097 43812
rect 44131 43809 44143 43843
rect 47412 43840 47440 43939
rect 47857 43843 47915 43849
rect 47857 43840 47869 43843
rect 47412 43812 47869 43840
rect 44085 43803 44143 43809
rect 47857 43809 47869 43812
rect 47903 43809 47915 43843
rect 47857 43803 47915 43809
rect 52546 43800 52552 43852
rect 52604 43800 52610 43852
rect 52730 43800 52736 43852
rect 52788 43800 52794 43852
rect 53929 43843 53987 43849
rect 53929 43809 53941 43843
rect 53975 43840 53987 43843
rect 66346 43840 66352 43852
rect 53975 43812 66352 43840
rect 53975 43809 53987 43812
rect 53929 43803 53987 43809
rect 44269 43775 44327 43781
rect 44269 43772 44281 43775
rect 43220 43744 44281 43772
rect 43220 43732 43226 43744
rect 44269 43741 44281 43744
rect 44315 43741 44327 43775
rect 44269 43735 44327 43741
rect 44910 43732 44916 43784
rect 44968 43772 44974 43784
rect 45097 43775 45155 43781
rect 45097 43772 45109 43775
rect 44968 43744 45109 43772
rect 44968 43732 44974 43744
rect 45097 43741 45109 43744
rect 45143 43741 45155 43775
rect 45097 43735 45155 43741
rect 45373 43775 45431 43781
rect 45373 43741 45385 43775
rect 45419 43772 45431 43775
rect 47394 43772 47400 43784
rect 45419 43744 47400 43772
rect 45419 43741 45431 43744
rect 45373 43735 45431 43741
rect 47394 43732 47400 43744
rect 47452 43732 47458 43784
rect 47486 43732 47492 43784
rect 47544 43732 47550 43784
rect 47673 43775 47731 43781
rect 47673 43741 47685 43775
rect 47719 43772 47731 43775
rect 47946 43772 47952 43784
rect 47719 43744 47952 43772
rect 47719 43741 47731 43744
rect 47673 43735 47731 43741
rect 47946 43732 47952 43744
rect 48004 43732 48010 43784
rect 41386 43676 42012 43704
rect 43625 43707 43683 43713
rect 43625 43673 43637 43707
rect 43671 43704 43683 43707
rect 44174 43704 44180 43716
rect 43671 43676 44180 43704
rect 43671 43673 43683 43676
rect 43625 43667 43683 43673
rect 44174 43664 44180 43676
rect 44232 43704 44238 43716
rect 44450 43704 44456 43716
rect 44232 43676 44456 43704
rect 44232 43664 44238 43676
rect 44450 43664 44456 43676
rect 44508 43664 44514 43716
rect 52917 43707 52975 43713
rect 52917 43673 52929 43707
rect 52963 43704 52975 43707
rect 53944 43704 53972 43803
rect 66346 43800 66352 43812
rect 66404 43800 66410 43852
rect 52963 43676 53972 43704
rect 52963 43673 52975 43676
rect 52917 43667 52975 43673
rect 35066 43636 35072 43648
rect 31812 43608 35072 43636
rect 31812 43596 31818 43608
rect 35066 43596 35072 43608
rect 35124 43596 35130 43648
rect 35250 43596 35256 43648
rect 35308 43596 35314 43648
rect 35526 43596 35532 43648
rect 35584 43596 35590 43648
rect 38562 43596 38568 43648
rect 38620 43596 38626 43648
rect 43806 43596 43812 43648
rect 43864 43596 43870 43648
rect 47029 43639 47087 43645
rect 47029 43605 47041 43639
rect 47075 43636 47087 43639
rect 47302 43636 47308 43648
rect 47075 43608 47308 43636
rect 47075 43605 47087 43608
rect 47029 43599 47087 43605
rect 47302 43596 47308 43608
rect 47360 43596 47366 43648
rect 48222 43596 48228 43648
rect 48280 43636 48286 43648
rect 48501 43639 48559 43645
rect 48501 43636 48513 43639
rect 48280 43608 48513 43636
rect 48280 43596 48286 43608
rect 48501 43605 48513 43608
rect 48547 43605 48559 43639
rect 48501 43599 48559 43605
rect 51902 43596 51908 43648
rect 51960 43636 51966 43648
rect 52273 43639 52331 43645
rect 52273 43636 52285 43639
rect 51960 43608 52285 43636
rect 51960 43596 51966 43608
rect 52273 43605 52285 43608
rect 52319 43605 52331 43639
rect 52273 43599 52331 43605
rect 53190 43596 53196 43648
rect 53248 43636 53254 43648
rect 53653 43639 53711 43645
rect 53653 43636 53665 43639
rect 53248 43608 53665 43636
rect 53248 43596 53254 43608
rect 53653 43605 53665 43608
rect 53699 43605 53711 43639
rect 53653 43599 53711 43605
rect 552 43546 66424 43568
rect 552 43494 1998 43546
rect 2050 43494 2062 43546
rect 2114 43494 2126 43546
rect 2178 43494 2190 43546
rect 2242 43494 2254 43546
rect 2306 43494 49998 43546
rect 50050 43494 50062 43546
rect 50114 43494 50126 43546
rect 50178 43494 50190 43546
rect 50242 43494 50254 43546
rect 50306 43494 66424 43546
rect 552 43472 66424 43494
rect 15378 43392 15384 43444
rect 15436 43432 15442 43444
rect 17405 43435 17463 43441
rect 17405 43432 17417 43435
rect 15436 43404 17417 43432
rect 15436 43392 15442 43404
rect 17405 43401 17417 43404
rect 17451 43401 17463 43435
rect 17405 43395 17463 43401
rect 17420 43364 17448 43395
rect 17494 43392 17500 43444
rect 17552 43392 17558 43444
rect 19518 43392 19524 43444
rect 19576 43432 19582 43444
rect 20441 43435 20499 43441
rect 20441 43432 20453 43435
rect 19576 43404 20453 43432
rect 19576 43392 19582 43404
rect 20441 43401 20453 43404
rect 20487 43432 20499 43435
rect 20530 43432 20536 43444
rect 20487 43404 20536 43432
rect 20487 43401 20499 43404
rect 20441 43395 20499 43401
rect 20530 43392 20536 43404
rect 20588 43392 20594 43444
rect 20640 43404 22508 43432
rect 18046 43364 18052 43376
rect 17420 43336 18052 43364
rect 18046 43324 18052 43336
rect 18104 43324 18110 43376
rect 20070 43324 20076 43376
rect 20128 43364 20134 43376
rect 20640 43364 20668 43404
rect 20128 43336 20668 43364
rect 22480 43364 22508 43404
rect 22554 43392 22560 43444
rect 22612 43392 22618 43444
rect 23382 43392 23388 43444
rect 23440 43432 23446 43444
rect 25593 43435 25651 43441
rect 25593 43432 25605 43435
rect 23440 43404 25605 43432
rect 23440 43392 23446 43404
rect 25593 43401 25605 43404
rect 25639 43432 25651 43435
rect 25774 43432 25780 43444
rect 25639 43404 25780 43432
rect 25639 43401 25651 43404
rect 25593 43395 25651 43401
rect 25774 43392 25780 43404
rect 25832 43392 25838 43444
rect 28810 43392 28816 43444
rect 28868 43392 28874 43444
rect 28902 43392 28908 43444
rect 28960 43432 28966 43444
rect 28960 43404 29408 43432
rect 28960 43392 28966 43404
rect 23290 43364 23296 43376
rect 22480 43336 23296 43364
rect 20128 43324 20134 43336
rect 23290 43324 23296 43336
rect 23348 43324 23354 43376
rect 25222 43324 25228 43376
rect 25280 43364 25286 43376
rect 25685 43367 25743 43373
rect 25685 43364 25697 43367
rect 25280 43336 25697 43364
rect 25280 43324 25286 43336
rect 25685 43333 25697 43336
rect 25731 43333 25743 43367
rect 26418 43364 26424 43376
rect 25685 43327 25743 43333
rect 26252 43336 26424 43364
rect 26252 43308 26280 43336
rect 26418 43324 26424 43336
rect 26476 43324 26482 43376
rect 27430 43364 27436 43376
rect 26712 43336 27436 43364
rect 13630 43256 13636 43308
rect 13688 43296 13694 43308
rect 15105 43299 15163 43305
rect 15105 43296 15117 43299
rect 13688 43268 15117 43296
rect 13688 43256 13694 43268
rect 15105 43265 15117 43268
rect 15151 43265 15163 43299
rect 15105 43259 15163 43265
rect 15657 43299 15715 43305
rect 15657 43265 15669 43299
rect 15703 43296 15715 43299
rect 15703 43268 18368 43296
rect 15703 43265 15715 43268
rect 15657 43259 15715 43265
rect 10686 43188 10692 43240
rect 10744 43188 10750 43240
rect 12098 43200 12434 43228
rect 10965 43163 11023 43169
rect 10965 43129 10977 43163
rect 11011 43160 11023 43163
rect 11238 43160 11244 43172
rect 11011 43132 11244 43160
rect 11011 43129 11023 43132
rect 10965 43123 11023 43129
rect 11238 43120 11244 43132
rect 11296 43120 11302 43172
rect 12406 43160 12434 43200
rect 15378 43188 15384 43240
rect 15436 43188 15442 43240
rect 18138 43188 18144 43240
rect 18196 43188 18202 43240
rect 18340 43228 18368 43268
rect 18414 43256 18420 43308
rect 18472 43256 18478 43308
rect 20809 43299 20867 43305
rect 20809 43296 20821 43299
rect 18708 43268 20821 43296
rect 18708 43237 18736 43268
rect 20809 43265 20821 43268
rect 20855 43265 20867 43299
rect 20809 43259 20867 43265
rect 23845 43299 23903 43305
rect 23845 43265 23857 43299
rect 23891 43296 23903 43299
rect 26234 43296 26240 43308
rect 23891 43268 26240 43296
rect 23891 43265 23903 43268
rect 23845 43259 23903 43265
rect 18693 43231 18751 43237
rect 18693 43228 18705 43231
rect 18340 43200 18705 43228
rect 18693 43197 18705 43200
rect 18739 43197 18751 43231
rect 18693 43191 18751 43197
rect 13814 43160 13820 43172
rect 12406 43132 13820 43160
rect 13814 43120 13820 43132
rect 13872 43160 13878 43172
rect 13872 43132 13938 43160
rect 13872 43120 13878 43132
rect 15930 43120 15936 43172
rect 15988 43120 15994 43172
rect 17678 43160 17684 43172
rect 17158 43132 17684 43160
rect 17678 43120 17684 43132
rect 17736 43120 17742 43172
rect 18966 43120 18972 43172
rect 19024 43120 19030 43172
rect 20346 43160 20352 43172
rect 20194 43132 20352 43160
rect 20346 43120 20352 43132
rect 20404 43120 20410 43172
rect 12437 43095 12495 43101
rect 12437 43061 12449 43095
rect 12483 43092 12495 43095
rect 12710 43092 12716 43104
rect 12483 43064 12716 43092
rect 12483 43061 12495 43064
rect 12437 43055 12495 43061
rect 12710 43052 12716 43064
rect 12768 43052 12774 43104
rect 12986 43052 12992 43104
rect 13044 43092 13050 43104
rect 13633 43095 13691 43101
rect 13633 43092 13645 43095
rect 13044 43064 13645 43092
rect 13044 43052 13050 43064
rect 13633 43061 13645 43064
rect 13679 43092 13691 43095
rect 13722 43092 13728 43104
rect 13679 43064 13728 43092
rect 13679 43061 13691 43064
rect 13633 43055 13691 43061
rect 13722 43052 13728 43064
rect 13780 43092 13786 43104
rect 15562 43092 15568 43104
rect 13780 43064 15568 43092
rect 13780 43052 13786 43064
rect 15562 43052 15568 43064
rect 15620 43052 15626 43104
rect 17770 43052 17776 43104
rect 17828 43052 17834 43104
rect 18233 43095 18291 43101
rect 18233 43061 18245 43095
rect 18279 43092 18291 43095
rect 19978 43092 19984 43104
rect 18279 43064 19984 43092
rect 18279 43061 18291 43064
rect 18233 43055 18291 43061
rect 19978 43052 19984 43064
rect 20036 43052 20042 43104
rect 20824 43092 20852 43259
rect 26234 43256 26240 43268
rect 26292 43256 26298 43308
rect 26329 43299 26387 43305
rect 26329 43265 26341 43299
rect 26375 43296 26387 43299
rect 26712 43296 26740 43336
rect 27430 43324 27436 43336
rect 27488 43324 27494 43376
rect 28074 43324 28080 43376
rect 28132 43364 28138 43376
rect 29273 43367 29331 43373
rect 29273 43364 29285 43367
rect 28132 43336 29285 43364
rect 28132 43324 28138 43336
rect 29273 43333 29285 43336
rect 29319 43333 29331 43367
rect 29380 43364 29408 43404
rect 29546 43392 29552 43444
rect 29604 43392 29610 43444
rect 29656 43404 33640 43432
rect 29656 43364 29684 43404
rect 29380 43336 29684 43364
rect 29273 43327 29331 43333
rect 26375 43268 26740 43296
rect 26789 43299 26847 43305
rect 26375 43265 26387 43268
rect 26329 43259 26387 43265
rect 26789 43265 26801 43299
rect 26835 43296 26847 43299
rect 27801 43299 27859 43305
rect 27801 43296 27813 43299
rect 26835 43268 27813 43296
rect 26835 43265 26847 43268
rect 26789 43259 26847 43265
rect 27801 43265 27813 43268
rect 27847 43296 27859 43299
rect 28261 43299 28319 43305
rect 28261 43296 28273 43299
rect 27847 43268 28273 43296
rect 27847 43265 27859 43268
rect 27801 43259 27859 43265
rect 28261 43265 28273 43268
rect 28307 43296 28319 43299
rect 28534 43296 28540 43308
rect 28307 43268 28540 43296
rect 28307 43265 28319 43268
rect 28261 43259 28319 43265
rect 22649 43231 22707 43237
rect 22649 43197 22661 43231
rect 22695 43228 22707 43231
rect 23474 43228 23480 43240
rect 22695 43200 23480 43228
rect 22695 43197 22707 43200
rect 22649 43191 22707 43197
rect 23474 43188 23480 43200
rect 23532 43188 23538 43240
rect 23658 43188 23664 43240
rect 23716 43188 23722 43240
rect 26050 43188 26056 43240
rect 26108 43228 26114 43240
rect 26344 43228 26372 43259
rect 28534 43256 28540 43268
rect 28592 43256 28598 43308
rect 29288 43296 29316 43327
rect 29914 43324 29920 43376
rect 29972 43364 29978 43376
rect 33612 43364 33640 43404
rect 34146 43392 34152 43444
rect 34204 43392 34210 43444
rect 34422 43392 34428 43444
rect 34480 43432 34486 43444
rect 34977 43435 35035 43441
rect 34977 43432 34989 43435
rect 34480 43404 34989 43432
rect 34480 43392 34486 43404
rect 34977 43401 34989 43404
rect 35023 43401 35035 43435
rect 34977 43395 35035 43401
rect 36354 43392 36360 43444
rect 36412 43392 36418 43444
rect 40773 43435 40831 43441
rect 40773 43401 40785 43435
rect 40819 43432 40831 43435
rect 40954 43432 40960 43444
rect 40819 43404 40960 43432
rect 40819 43401 40831 43404
rect 40773 43395 40831 43401
rect 40954 43392 40960 43404
rect 41012 43392 41018 43444
rect 42334 43392 42340 43444
rect 42392 43432 42398 43444
rect 43533 43435 43591 43441
rect 43533 43432 43545 43435
rect 42392 43404 43545 43432
rect 42392 43392 42398 43404
rect 43533 43401 43545 43404
rect 43579 43401 43591 43435
rect 43533 43395 43591 43401
rect 43806 43392 43812 43444
rect 43864 43432 43870 43444
rect 43864 43404 44128 43432
rect 43864 43392 43870 43404
rect 35434 43364 35440 43376
rect 29972 43336 31892 43364
rect 33612 43336 35440 43364
rect 29972 43324 29978 43336
rect 30101 43299 30159 43305
rect 30101 43296 30113 43299
rect 29288 43268 30113 43296
rect 30101 43265 30113 43268
rect 30147 43265 30159 43299
rect 30101 43259 30159 43265
rect 30208 43268 31432 43296
rect 26108 43200 26372 43228
rect 26973 43231 27031 43237
rect 26108 43188 26114 43200
rect 26973 43197 26985 43231
rect 27019 43228 27031 43231
rect 28350 43228 28356 43240
rect 27019 43200 28356 43228
rect 27019 43197 27031 43200
rect 26973 43191 27031 43197
rect 28350 43188 28356 43200
rect 28408 43188 28414 43240
rect 28445 43231 28503 43237
rect 28445 43197 28457 43231
rect 28491 43228 28503 43231
rect 29914 43228 29920 43240
rect 28491 43200 29920 43228
rect 28491 43197 28503 43200
rect 28445 43191 28503 43197
rect 29914 43188 29920 43200
rect 29972 43188 29978 43240
rect 21085 43163 21143 43169
rect 21085 43129 21097 43163
rect 21131 43160 21143 43163
rect 21174 43160 21180 43172
rect 21131 43132 21180 43160
rect 21131 43129 21143 43132
rect 21085 43123 21143 43129
rect 21174 43120 21180 43132
rect 21232 43120 21238 43172
rect 21634 43120 21640 43172
rect 21692 43120 21698 43172
rect 24121 43163 24179 43169
rect 24121 43129 24133 43163
rect 24167 43160 24179 43163
rect 24210 43160 24216 43172
rect 24167 43132 24216 43160
rect 24167 43129 24179 43132
rect 24121 43123 24179 43129
rect 24210 43120 24216 43132
rect 24268 43120 24274 43172
rect 24854 43120 24860 43172
rect 24912 43120 24918 43172
rect 26881 43163 26939 43169
rect 26881 43160 26893 43163
rect 26068 43132 26893 43160
rect 22002 43092 22008 43104
rect 20824 43064 22008 43092
rect 22002 43052 22008 43064
rect 22060 43052 22066 43104
rect 22830 43052 22836 43104
rect 22888 43052 22894 43104
rect 23014 43052 23020 43104
rect 23072 43052 23078 43104
rect 25406 43052 25412 43104
rect 25464 43092 25470 43104
rect 25866 43092 25872 43104
rect 25464 43064 25872 43092
rect 25464 43052 25470 43064
rect 25866 43052 25872 43064
rect 25924 43092 25930 43104
rect 26068 43101 26096 43132
rect 26881 43129 26893 43132
rect 26927 43129 26939 43163
rect 26881 43123 26939 43129
rect 27522 43120 27528 43172
rect 27580 43160 27586 43172
rect 28902 43160 28908 43172
rect 27580 43132 28908 43160
rect 27580 43120 27586 43132
rect 28902 43120 28908 43132
rect 28960 43120 28966 43172
rect 29089 43163 29147 43169
rect 29089 43129 29101 43163
rect 29135 43160 29147 43163
rect 30208 43160 30236 43268
rect 30282 43188 30288 43240
rect 30340 43228 30346 43240
rect 31297 43231 31355 43237
rect 31297 43228 31309 43231
rect 30340 43200 31309 43228
rect 30340 43188 30346 43200
rect 31297 43197 31309 43200
rect 31343 43197 31355 43231
rect 31404 43228 31432 43268
rect 31754 43256 31760 43308
rect 31812 43256 31818 43308
rect 31864 43296 31892 43336
rect 35434 43324 35440 43336
rect 35492 43324 35498 43376
rect 39390 43324 39396 43376
rect 39448 43364 39454 43376
rect 39448 43336 41184 43364
rect 39448 43324 39454 43336
rect 33318 43296 33324 43308
rect 31864 43268 33324 43296
rect 33318 43256 33324 43268
rect 33376 43256 33382 43308
rect 34793 43299 34851 43305
rect 34793 43296 34805 43299
rect 34440 43268 34805 43296
rect 33873 43231 33931 43237
rect 31404 43200 31754 43228
rect 31297 43191 31355 43197
rect 29135 43132 30236 43160
rect 30469 43163 30527 43169
rect 29135 43129 29147 43132
rect 29089 43123 29147 43129
rect 30469 43129 30481 43163
rect 30515 43160 30527 43163
rect 31202 43160 31208 43172
rect 30515 43132 31208 43160
rect 30515 43129 30527 43132
rect 30469 43123 30527 43129
rect 26053 43095 26111 43101
rect 26053 43092 26065 43095
rect 25924 43064 26065 43092
rect 25924 43052 25930 43064
rect 26053 43061 26065 43064
rect 26099 43061 26111 43095
rect 26053 43055 26111 43061
rect 26145 43095 26203 43101
rect 26145 43061 26157 43095
rect 26191 43092 26203 43095
rect 26234 43092 26240 43104
rect 26191 43064 26240 43092
rect 26191 43061 26203 43064
rect 26145 43055 26203 43061
rect 26234 43052 26240 43064
rect 26292 43052 26298 43104
rect 27338 43052 27344 43104
rect 27396 43052 27402 43104
rect 27430 43052 27436 43104
rect 27488 43092 27494 43104
rect 29104 43092 29132 43123
rect 31202 43120 31208 43132
rect 31260 43120 31266 43172
rect 27488 43064 29132 43092
rect 27488 43052 27494 43064
rect 30006 43052 30012 43104
rect 30064 43052 30070 43104
rect 30558 43052 30564 43104
rect 30616 43052 30622 43104
rect 31294 43052 31300 43104
rect 31352 43092 31358 43104
rect 31389 43095 31447 43101
rect 31389 43092 31401 43095
rect 31352 43064 31401 43092
rect 31352 43052 31358 43064
rect 31389 43061 31401 43064
rect 31435 43061 31447 43095
rect 31726 43092 31754 43200
rect 33873 43197 33885 43231
rect 33919 43228 33931 43231
rect 34440 43228 34468 43268
rect 34793 43265 34805 43268
rect 34839 43296 34851 43299
rect 35158 43296 35164 43308
rect 34839 43268 35164 43296
rect 34839 43265 34851 43268
rect 34793 43259 34851 43265
rect 35158 43256 35164 43268
rect 35216 43256 35222 43308
rect 35529 43299 35587 43305
rect 35529 43265 35541 43299
rect 35575 43265 35587 43299
rect 35529 43259 35587 43265
rect 33919 43200 34468 43228
rect 33919 43197 33931 43200
rect 33873 43191 33931 43197
rect 34514 43188 34520 43240
rect 34572 43188 34578 43240
rect 35250 43188 35256 43240
rect 35308 43228 35314 43240
rect 35345 43231 35403 43237
rect 35345 43228 35357 43231
rect 35308 43200 35357 43228
rect 35308 43188 35314 43200
rect 35345 43197 35357 43200
rect 35391 43197 35403 43231
rect 35345 43191 35403 43197
rect 32030 43120 32036 43172
rect 32088 43120 32094 43172
rect 32490 43120 32496 43172
rect 32548 43120 32554 43172
rect 33689 43163 33747 43169
rect 33689 43160 33701 43163
rect 33336 43132 33701 43160
rect 33336 43092 33364 43132
rect 33689 43129 33701 43132
rect 33735 43129 33747 43163
rect 33689 43123 33747 43129
rect 34422 43120 34428 43172
rect 34480 43160 34486 43172
rect 35437 43163 35495 43169
rect 35437 43160 35449 43163
rect 34480 43132 35449 43160
rect 34480 43120 34486 43132
rect 35437 43129 35449 43132
rect 35483 43129 35495 43163
rect 35437 43123 35495 43129
rect 31726 43064 33364 43092
rect 33505 43095 33563 43101
rect 31389 43055 31447 43061
rect 33505 43061 33517 43095
rect 33551 43092 33563 43095
rect 34440 43092 34468 43120
rect 33551 43064 34468 43092
rect 34609 43095 34667 43101
rect 33551 43061 33563 43064
rect 33505 43055 33563 43061
rect 34609 43061 34621 43095
rect 34655 43092 34667 43095
rect 34790 43092 34796 43104
rect 34655 43064 34796 43092
rect 34655 43061 34667 43064
rect 34609 43055 34667 43061
rect 34790 43052 34796 43064
rect 34848 43052 34854 43104
rect 35342 43052 35348 43104
rect 35400 43092 35406 43104
rect 35544 43092 35572 43259
rect 38286 43256 38292 43308
rect 38344 43296 38350 43308
rect 38749 43299 38807 43305
rect 38749 43296 38761 43299
rect 38344 43268 38761 43296
rect 38344 43256 38350 43268
rect 38749 43265 38761 43268
rect 38795 43265 38807 43299
rect 38749 43259 38807 43265
rect 40126 43256 40132 43308
rect 40184 43296 40190 43308
rect 40497 43299 40555 43305
rect 40497 43296 40509 43299
rect 40184 43268 40509 43296
rect 40184 43256 40190 43268
rect 40497 43265 40509 43268
rect 40543 43265 40555 43299
rect 40497 43259 40555 43265
rect 41156 43296 41184 43336
rect 41230 43324 41236 43376
rect 41288 43364 41294 43376
rect 41288 43336 41736 43364
rect 41288 43324 41294 43336
rect 41156 43268 41368 43296
rect 38105 43231 38163 43237
rect 38105 43197 38117 43231
rect 38151 43197 38163 43231
rect 38105 43191 38163 43197
rect 37734 43160 37740 43172
rect 37398 43132 37740 43160
rect 37734 43120 37740 43132
rect 37792 43120 37798 43172
rect 37829 43163 37887 43169
rect 37829 43129 37841 43163
rect 37875 43129 37887 43163
rect 37829 43123 37887 43129
rect 35400 43064 35572 43092
rect 37844 43092 37872 43123
rect 37918 43120 37924 43172
rect 37976 43160 37982 43172
rect 38120 43160 38148 43191
rect 38562 43188 38568 43240
rect 38620 43188 38626 43240
rect 40310 43188 40316 43240
rect 40368 43188 40374 43240
rect 41156 43237 41184 43268
rect 41141 43231 41199 43237
rect 41141 43197 41153 43231
rect 41187 43197 41199 43231
rect 41340 43228 41368 43268
rect 41414 43256 41420 43308
rect 41472 43256 41478 43308
rect 41708 43305 41736 43336
rect 43346 43324 43352 43376
rect 43404 43364 43410 43376
rect 43441 43367 43499 43373
rect 43441 43364 43453 43367
rect 43404 43336 43453 43364
rect 43404 43324 43410 43336
rect 43441 43333 43453 43336
rect 43487 43364 43499 43367
rect 43487 43336 44036 43364
rect 43487 43333 43499 43336
rect 43441 43327 43499 43333
rect 44008 43308 44036 43336
rect 44100 43308 44128 43404
rect 47486 43392 47492 43444
rect 47544 43432 47550 43444
rect 48777 43435 48835 43441
rect 48777 43432 48789 43435
rect 47544 43404 48789 43432
rect 47544 43392 47550 43404
rect 48777 43401 48789 43404
rect 48823 43401 48835 43435
rect 48777 43395 48835 43401
rect 49510 43392 49516 43444
rect 49568 43432 49574 43444
rect 49568 43404 51948 43432
rect 49568 43392 49574 43404
rect 51920 43364 51948 43404
rect 52546 43392 52552 43444
rect 52604 43432 52610 43444
rect 53929 43435 53987 43441
rect 53929 43432 53941 43435
rect 52604 43404 53941 43432
rect 52604 43392 52610 43404
rect 53929 43401 53941 43404
rect 53975 43432 53987 43435
rect 53975 43404 55214 43432
rect 53975 43401 53987 43404
rect 53929 43395 53987 43401
rect 51920 43336 53328 43364
rect 41693 43299 41751 43305
rect 41693 43265 41705 43299
rect 41739 43296 41751 43299
rect 41739 43268 43300 43296
rect 41739 43265 41751 43268
rect 41693 43259 41751 43265
rect 41340 43200 41414 43228
rect 41141 43191 41199 43197
rect 37976 43132 38148 43160
rect 37976 43120 37982 43132
rect 38838 43120 38844 43172
rect 38896 43160 38902 43172
rect 39390 43160 39396 43172
rect 38896 43132 39396 43160
rect 38896 43120 38902 43132
rect 39390 43120 39396 43132
rect 39448 43120 39454 43172
rect 41386 43160 41414 43200
rect 43070 43188 43076 43240
rect 43128 43188 43134 43240
rect 43272 43228 43300 43268
rect 43990 43256 43996 43308
rect 44048 43256 44054 43308
rect 44082 43256 44088 43308
rect 44140 43256 44146 43308
rect 45370 43256 45376 43308
rect 45428 43256 45434 43308
rect 45922 43256 45928 43308
rect 45980 43296 45986 43308
rect 46842 43296 46848 43308
rect 45980 43268 46848 43296
rect 45980 43256 45986 43268
rect 46842 43256 46848 43268
rect 46900 43256 46906 43308
rect 47302 43256 47308 43308
rect 47360 43256 47366 43308
rect 50617 43299 50675 43305
rect 50617 43265 50629 43299
rect 50663 43296 50675 43299
rect 51258 43296 51264 43308
rect 50663 43268 51264 43296
rect 50663 43265 50675 43268
rect 50617 43259 50675 43265
rect 51258 43256 51264 43268
rect 51316 43256 51322 43308
rect 52365 43299 52423 43305
rect 52365 43265 52377 43299
rect 52411 43296 52423 43299
rect 52546 43296 52552 43308
rect 52411 43268 52552 43296
rect 52411 43265 52423 43268
rect 52365 43259 52423 43265
rect 52546 43256 52552 43268
rect 52604 43296 52610 43308
rect 53009 43299 53067 43305
rect 53009 43296 53021 43299
rect 52604 43268 53021 43296
rect 52604 43256 52610 43268
rect 53009 43265 53021 43268
rect 53055 43265 53067 43299
rect 53009 43259 53067 43265
rect 44818 43228 44824 43240
rect 43272 43200 44824 43228
rect 44818 43188 44824 43200
rect 44876 43228 44882 43240
rect 45097 43231 45155 43237
rect 45097 43228 45109 43231
rect 44876 43200 45109 43228
rect 44876 43188 44882 43200
rect 45097 43197 45109 43200
rect 45143 43197 45155 43231
rect 45097 43191 45155 43197
rect 46934 43188 46940 43240
rect 46992 43228 46998 43240
rect 53300 43237 53328 43336
rect 47029 43231 47087 43237
rect 47029 43228 47041 43231
rect 46992 43200 47041 43228
rect 46992 43188 46998 43200
rect 47029 43197 47041 43200
rect 47075 43197 47087 43231
rect 47029 43191 47087 43197
rect 53285 43231 53343 43237
rect 53285 43197 53297 43231
rect 53331 43197 53343 43231
rect 53285 43191 53343 43197
rect 53834 43188 53840 43240
rect 53892 43188 53898 43240
rect 41386 43132 41920 43160
rect 38197 43095 38255 43101
rect 38197 43092 38209 43095
rect 37844 43064 38209 43092
rect 35400 43052 35406 43064
rect 38197 43061 38209 43064
rect 38243 43061 38255 43095
rect 38197 43055 38255 43061
rect 38378 43052 38384 43104
rect 38436 43092 38442 43104
rect 38657 43095 38715 43101
rect 38657 43092 38669 43095
rect 38436 43064 38669 43092
rect 38436 43052 38442 43064
rect 38657 43061 38669 43064
rect 38703 43061 38715 43095
rect 38657 43055 38715 43061
rect 39298 43052 39304 43104
rect 39356 43092 39362 43104
rect 39485 43095 39543 43101
rect 39485 43092 39497 43095
rect 39356 43064 39497 43092
rect 39356 43052 39362 43064
rect 39485 43061 39497 43064
rect 39531 43061 39543 43095
rect 39485 43055 39543 43061
rect 39574 43052 39580 43104
rect 39632 43092 39638 43104
rect 39945 43095 40003 43101
rect 39945 43092 39957 43095
rect 39632 43064 39957 43092
rect 39632 43052 39638 43064
rect 39945 43061 39957 43064
rect 39991 43061 40003 43095
rect 39945 43055 40003 43061
rect 40402 43052 40408 43104
rect 40460 43052 40466 43104
rect 41233 43095 41291 43101
rect 41233 43061 41245 43095
rect 41279 43092 41291 43095
rect 41782 43092 41788 43104
rect 41279 43064 41788 43092
rect 41279 43061 41291 43064
rect 41233 43055 41291 43061
rect 41782 43052 41788 43064
rect 41840 43052 41846 43104
rect 41892 43092 41920 43132
rect 41966 43120 41972 43172
rect 42024 43120 42030 43172
rect 43901 43163 43959 43169
rect 43901 43160 43913 43163
rect 43272 43132 43913 43160
rect 43272 43092 43300 43132
rect 43901 43129 43913 43132
rect 43947 43129 43959 43163
rect 46658 43160 46664 43172
rect 46598 43132 46664 43160
rect 43901 43123 43959 43129
rect 46658 43120 46664 43132
rect 46716 43160 46722 43172
rect 48958 43160 48964 43172
rect 46716 43132 47716 43160
rect 48530 43132 48964 43160
rect 46716 43120 46722 43132
rect 41892 43064 43300 43092
rect 47688 43092 47716 43132
rect 48608 43092 48636 43132
rect 48958 43120 48964 43132
rect 49016 43120 49022 43172
rect 50893 43163 50951 43169
rect 50893 43129 50905 43163
rect 50939 43160 50951 43163
rect 53190 43160 53196 43172
rect 50939 43132 51074 43160
rect 52118 43132 53196 43160
rect 50939 43129 50951 43132
rect 50893 43123 50951 43129
rect 47688 43064 48636 43092
rect 51046 43092 51074 43132
rect 53190 43120 53196 43132
rect 53248 43120 53254 43172
rect 51534 43092 51540 43104
rect 51046 43064 51540 43092
rect 51534 43052 51540 43064
rect 51592 43052 51598 43104
rect 52454 43052 52460 43104
rect 52512 43052 52518 43104
rect 53374 43052 53380 43104
rect 53432 43052 53438 43104
rect 55186 43092 55214 43404
rect 60642 43092 60648 43104
rect 55186 43064 60648 43092
rect 60642 43052 60648 43064
rect 60700 43052 60706 43104
rect 552 43002 66424 43024
rect 552 42950 2918 43002
rect 2970 42950 2982 43002
rect 3034 42950 3046 43002
rect 3098 42950 3110 43002
rect 3162 42950 3174 43002
rect 3226 42950 50918 43002
rect 50970 42950 50982 43002
rect 51034 42950 51046 43002
rect 51098 42950 51110 43002
rect 51162 42950 51174 43002
rect 51226 42950 66424 43002
rect 552 42928 66424 42950
rect 11238 42848 11244 42900
rect 11296 42888 11302 42900
rect 11333 42891 11391 42897
rect 11333 42888 11345 42891
rect 11296 42860 11345 42888
rect 11296 42848 11302 42860
rect 11333 42857 11345 42860
rect 11379 42857 11391 42891
rect 11333 42851 11391 42857
rect 11698 42848 11704 42900
rect 11756 42848 11762 42900
rect 14553 42891 14611 42897
rect 14553 42857 14565 42891
rect 14599 42888 14611 42891
rect 14642 42888 14648 42900
rect 14599 42860 14648 42888
rect 14599 42857 14611 42860
rect 14553 42851 14611 42857
rect 14642 42848 14648 42860
rect 14700 42848 14706 42900
rect 15194 42848 15200 42900
rect 15252 42848 15258 42900
rect 16850 42848 16856 42900
rect 16908 42848 16914 42900
rect 17678 42848 17684 42900
rect 17736 42888 17742 42900
rect 17736 42860 19196 42888
rect 17736 42848 17742 42860
rect 13814 42780 13820 42832
rect 13872 42780 13878 42832
rect 15562 42780 15568 42832
rect 15620 42780 15626 42832
rect 15657 42823 15715 42829
rect 15657 42789 15669 42823
rect 15703 42820 15715 42823
rect 15703 42792 16436 42820
rect 15703 42789 15715 42792
rect 15657 42783 15715 42789
rect 11793 42755 11851 42761
rect 11793 42721 11805 42755
rect 11839 42752 11851 42755
rect 12710 42752 12716 42764
rect 11839 42724 12716 42752
rect 11839 42721 11851 42724
rect 11793 42715 11851 42721
rect 12710 42712 12716 42724
rect 12768 42712 12774 42764
rect 15105 42755 15163 42761
rect 15105 42721 15117 42755
rect 15151 42752 15163 42755
rect 15672 42752 15700 42783
rect 15151 42724 15700 42752
rect 15151 42721 15163 42724
rect 15105 42715 15163 42721
rect 15838 42712 15844 42764
rect 15896 42752 15902 42764
rect 16117 42755 16175 42761
rect 16117 42752 16129 42755
rect 15896 42724 16129 42752
rect 15896 42712 15902 42724
rect 16117 42721 16129 42724
rect 16163 42721 16175 42755
rect 16408 42752 16436 42792
rect 16482 42780 16488 42832
rect 16540 42820 16546 42832
rect 17126 42820 17132 42832
rect 16540 42792 17132 42820
rect 16540 42780 16546 42792
rect 17126 42780 17132 42792
rect 17184 42780 17190 42832
rect 17770 42780 17776 42832
rect 17828 42820 17834 42832
rect 17865 42823 17923 42829
rect 17865 42820 17877 42823
rect 17828 42792 17877 42820
rect 17828 42780 17834 42792
rect 17865 42789 17877 42792
rect 17911 42789 17923 42823
rect 19168 42820 19196 42860
rect 19334 42848 19340 42900
rect 19392 42848 19398 42900
rect 19978 42848 19984 42900
rect 20036 42888 20042 42900
rect 20073 42891 20131 42897
rect 20073 42888 20085 42891
rect 20036 42860 20085 42888
rect 20036 42848 20042 42860
rect 20073 42857 20085 42860
rect 20119 42857 20131 42891
rect 20073 42851 20131 42857
rect 20438 42848 20444 42900
rect 20496 42848 20502 42900
rect 20530 42848 20536 42900
rect 20588 42848 20594 42900
rect 21913 42891 21971 42897
rect 21913 42857 21925 42891
rect 21959 42888 21971 42891
rect 21959 42860 23152 42888
rect 21959 42857 21971 42860
rect 21913 42851 21971 42857
rect 19889 42823 19947 42829
rect 19090 42792 19380 42820
rect 17865 42783 17923 42789
rect 16408 42724 17264 42752
rect 16117 42715 16175 42721
rect 9490 42644 9496 42696
rect 9548 42644 9554 42696
rect 11977 42687 12035 42693
rect 11977 42653 11989 42687
rect 12023 42684 12035 42687
rect 12618 42684 12624 42696
rect 12023 42656 12624 42684
rect 12023 42653 12035 42656
rect 11977 42647 12035 42653
rect 12618 42644 12624 42656
rect 12676 42644 12682 42696
rect 12802 42644 12808 42696
rect 12860 42644 12866 42696
rect 13081 42687 13139 42693
rect 13081 42653 13093 42687
rect 13127 42684 13139 42687
rect 14458 42684 14464 42696
rect 13127 42656 14464 42684
rect 13127 42653 13139 42656
rect 13081 42647 13139 42653
rect 14458 42644 14464 42656
rect 14516 42644 14522 42696
rect 15749 42687 15807 42693
rect 15749 42653 15761 42687
rect 15795 42684 15807 42687
rect 16666 42684 16672 42696
rect 15795 42656 16672 42684
rect 15795 42653 15807 42656
rect 15749 42647 15807 42653
rect 8938 42508 8944 42560
rect 8996 42508 9002 42560
rect 13170 42508 13176 42560
rect 13228 42548 13234 42560
rect 13538 42548 13544 42560
rect 13228 42520 13544 42548
rect 13228 42508 13234 42520
rect 13538 42508 13544 42520
rect 13596 42548 13602 42560
rect 15764 42548 15792 42647
rect 16666 42644 16672 42656
rect 16724 42644 16730 42696
rect 16942 42644 16948 42696
rect 17000 42644 17006 42696
rect 17126 42644 17132 42696
rect 17184 42644 17190 42696
rect 17236 42684 17264 42724
rect 17310 42712 17316 42764
rect 17368 42712 17374 42764
rect 17586 42712 17592 42764
rect 17644 42712 17650 42764
rect 19352 42752 19380 42792
rect 19889 42789 19901 42823
rect 19935 42820 19947 42823
rect 20456 42820 20484 42848
rect 19935 42792 20484 42820
rect 22373 42823 22431 42829
rect 19935 42789 19947 42792
rect 19889 42783 19947 42789
rect 22373 42789 22385 42823
rect 22419 42820 22431 42823
rect 22646 42820 22652 42832
rect 22419 42792 22652 42820
rect 22419 42789 22431 42792
rect 22373 42783 22431 42789
rect 22646 42780 22652 42792
rect 22704 42780 22710 42832
rect 22830 42780 22836 42832
rect 22888 42780 22894 42832
rect 23124 42829 23152 42860
rect 23474 42848 23480 42900
rect 23532 42888 23538 42900
rect 24946 42888 24952 42900
rect 23532 42860 24952 42888
rect 23532 42848 23538 42860
rect 24946 42848 24952 42860
rect 25004 42848 25010 42900
rect 25774 42848 25780 42900
rect 25832 42848 25838 42900
rect 25869 42891 25927 42897
rect 25869 42857 25881 42891
rect 25915 42888 25927 42891
rect 25958 42888 25964 42900
rect 25915 42860 25964 42888
rect 25915 42857 25927 42860
rect 25869 42851 25927 42857
rect 25958 42848 25964 42860
rect 26016 42848 26022 42900
rect 26234 42848 26240 42900
rect 26292 42848 26298 42900
rect 26326 42848 26332 42900
rect 26384 42888 26390 42900
rect 26421 42891 26479 42897
rect 26421 42888 26433 42891
rect 26384 42860 26433 42888
rect 26384 42848 26390 42860
rect 26421 42857 26433 42860
rect 26467 42857 26479 42891
rect 26421 42851 26479 42857
rect 27157 42891 27215 42897
rect 27157 42857 27169 42891
rect 27203 42888 27215 42891
rect 27338 42888 27344 42900
rect 27203 42860 27344 42888
rect 27203 42857 27215 42860
rect 27157 42851 27215 42857
rect 27338 42848 27344 42860
rect 27396 42848 27402 42900
rect 27982 42848 27988 42900
rect 28040 42848 28046 42900
rect 29917 42891 29975 42897
rect 29917 42857 29929 42891
rect 29963 42888 29975 42891
rect 30006 42888 30012 42900
rect 29963 42860 30012 42888
rect 29963 42857 29975 42860
rect 29917 42851 29975 42857
rect 30006 42848 30012 42860
rect 30064 42848 30070 42900
rect 30558 42848 30564 42900
rect 30616 42888 30622 42900
rect 31754 42888 31760 42900
rect 30616 42860 31760 42888
rect 30616 42848 30622 42860
rect 31754 42848 31760 42860
rect 31812 42888 31818 42900
rect 32490 42888 32496 42900
rect 31812 42860 32496 42888
rect 31812 42848 31818 42860
rect 32490 42848 32496 42860
rect 32548 42848 32554 42900
rect 32582 42848 32588 42900
rect 32640 42888 32646 42900
rect 32677 42891 32735 42897
rect 32677 42888 32689 42891
rect 32640 42860 32689 42888
rect 32640 42848 32646 42860
rect 32677 42857 32689 42860
rect 32723 42857 32735 42891
rect 32677 42851 32735 42857
rect 33042 42848 33048 42900
rect 33100 42848 33106 42900
rect 34330 42848 34336 42900
rect 34388 42848 34394 42900
rect 34790 42848 34796 42900
rect 34848 42848 34854 42900
rect 36081 42891 36139 42897
rect 36081 42857 36093 42891
rect 36127 42888 36139 42891
rect 36722 42888 36728 42900
rect 36127 42860 36728 42888
rect 36127 42857 36139 42860
rect 36081 42851 36139 42857
rect 36722 42848 36728 42860
rect 36780 42848 36786 42900
rect 39482 42848 39488 42900
rect 39540 42848 39546 42900
rect 40129 42891 40187 42897
rect 40129 42857 40141 42891
rect 40175 42857 40187 42891
rect 40129 42851 40187 42857
rect 23109 42823 23167 42829
rect 23109 42789 23121 42823
rect 23155 42789 23167 42823
rect 24854 42820 24860 42832
rect 24334 42792 24860 42820
rect 23109 42783 23167 42789
rect 24854 42780 24860 42792
rect 24912 42780 24918 42832
rect 27065 42823 27123 42829
rect 26160 42792 27016 42820
rect 20346 42752 20352 42764
rect 19352 42724 20352 42752
rect 20346 42712 20352 42724
rect 20404 42712 20410 42764
rect 22281 42755 22339 42761
rect 22281 42721 22293 42755
rect 22327 42752 22339 42755
rect 22554 42752 22560 42764
rect 22327 42724 22560 42752
rect 22327 42721 22339 42724
rect 22281 42715 22339 42721
rect 22554 42712 22560 42724
rect 22612 42712 22618 42764
rect 22848 42752 22876 42780
rect 25038 42752 25044 42764
rect 22756 42724 22876 42752
rect 24596 42724 25044 42752
rect 17236 42656 19334 42684
rect 16022 42576 16028 42628
rect 16080 42616 16086 42628
rect 19306 42616 19334 42656
rect 20530 42644 20536 42696
rect 20588 42684 20594 42696
rect 20625 42687 20683 42693
rect 20625 42684 20637 42687
rect 20588 42656 20637 42684
rect 20588 42644 20594 42656
rect 20625 42653 20637 42656
rect 20671 42653 20683 42687
rect 20625 42647 20683 42653
rect 21358 42644 21364 42696
rect 21416 42644 21422 42696
rect 22097 42687 22155 42693
rect 22097 42653 22109 42687
rect 22143 42684 22155 42687
rect 22756 42684 22784 42724
rect 24596 42693 24624 42724
rect 25038 42712 25044 42724
rect 25096 42712 25102 42764
rect 26050 42752 26056 42764
rect 25332 42724 26056 42752
rect 22143 42656 22784 42684
rect 22833 42687 22891 42693
rect 22143 42653 22155 42656
rect 22097 42647 22155 42653
rect 22833 42653 22845 42687
rect 22879 42653 22891 42687
rect 22833 42647 22891 42653
rect 24581 42687 24639 42693
rect 24581 42653 24593 42687
rect 24627 42653 24639 42687
rect 24581 42647 24639 42653
rect 21266 42616 21272 42628
rect 16080 42588 16712 42616
rect 19306 42588 21272 42616
rect 16080 42576 16086 42588
rect 13596 42520 15792 42548
rect 13596 42508 13602 42520
rect 16298 42508 16304 42560
rect 16356 42508 16362 42560
rect 16390 42508 16396 42560
rect 16448 42548 16454 42560
rect 16485 42551 16543 42557
rect 16485 42548 16497 42551
rect 16448 42520 16497 42548
rect 16448 42508 16454 42520
rect 16485 42517 16497 42520
rect 16531 42517 16543 42551
rect 16684 42548 16712 42588
rect 21266 42576 21272 42588
rect 21324 42576 21330 42628
rect 22186 42576 22192 42628
rect 22244 42616 22250 42628
rect 22848 42616 22876 42647
rect 24670 42644 24676 42696
rect 24728 42684 24734 42696
rect 24728 42656 25084 42684
rect 24728 42644 24734 42656
rect 24946 42616 24952 42628
rect 22244 42588 22876 42616
rect 24136 42588 24952 42616
rect 22244 42576 22250 42588
rect 17586 42548 17592 42560
rect 16684 42520 17592 42548
rect 16485 42511 16543 42517
rect 17586 42508 17592 42520
rect 17644 42548 17650 42560
rect 20162 42548 20168 42560
rect 17644 42520 20168 42548
rect 17644 42508 17650 42520
rect 20162 42508 20168 42520
rect 20220 42508 20226 42560
rect 20530 42508 20536 42560
rect 20588 42548 20594 42560
rect 22370 42548 22376 42560
rect 20588 42520 22376 42548
rect 20588 42508 20594 42520
rect 22370 42508 22376 42520
rect 22428 42508 22434 42560
rect 22554 42508 22560 42560
rect 22612 42548 22618 42560
rect 22741 42551 22799 42557
rect 22741 42548 22753 42551
rect 22612 42520 22753 42548
rect 22612 42508 22618 42520
rect 22741 42517 22753 42520
rect 22787 42517 22799 42551
rect 22741 42511 22799 42517
rect 22830 42508 22836 42560
rect 22888 42548 22894 42560
rect 24136 42548 24164 42588
rect 24946 42576 24952 42588
rect 25004 42576 25010 42628
rect 22888 42520 24164 42548
rect 22888 42508 22894 42520
rect 24210 42508 24216 42560
rect 24268 42548 24274 42560
rect 24673 42551 24731 42557
rect 24673 42548 24685 42551
rect 24268 42520 24685 42548
rect 24268 42508 24274 42520
rect 24673 42517 24685 42520
rect 24719 42517 24731 42551
rect 25056 42548 25084 42656
rect 25130 42644 25136 42696
rect 25188 42644 25194 42696
rect 25222 42644 25228 42696
rect 25280 42684 25286 42696
rect 25332 42693 25360 42724
rect 26050 42712 26056 42724
rect 26108 42712 26114 42764
rect 25317 42687 25375 42693
rect 25317 42684 25329 42687
rect 25280 42656 25329 42684
rect 25280 42644 25286 42656
rect 25317 42653 25329 42656
rect 25363 42653 25375 42687
rect 25317 42647 25375 42653
rect 25682 42644 25688 42696
rect 25740 42684 25746 42696
rect 26160 42684 26188 42792
rect 26510 42712 26516 42764
rect 26568 42752 26574 42764
rect 26605 42755 26663 42761
rect 26605 42752 26617 42755
rect 26568 42724 26617 42752
rect 26568 42712 26574 42724
rect 26605 42721 26617 42724
rect 26651 42721 26663 42755
rect 26988 42752 27016 42792
rect 27065 42789 27077 42823
rect 27111 42820 27123 42823
rect 29089 42823 29147 42829
rect 29089 42820 29101 42823
rect 27111 42792 29101 42820
rect 27111 42789 27123 42792
rect 27065 42783 27123 42789
rect 29089 42789 29101 42792
rect 29135 42789 29147 42823
rect 29089 42783 29147 42789
rect 30285 42823 30343 42829
rect 30285 42789 30297 42823
rect 30331 42820 30343 42823
rect 30650 42820 30656 42832
rect 30331 42792 30656 42820
rect 30331 42789 30343 42792
rect 30285 42783 30343 42789
rect 30650 42780 30656 42792
rect 30708 42780 30714 42832
rect 36170 42780 36176 42832
rect 36228 42780 36234 42832
rect 36354 42780 36360 42832
rect 36412 42820 36418 42832
rect 37001 42823 37059 42829
rect 37001 42820 37013 42823
rect 36412 42792 37013 42820
rect 36412 42780 36418 42792
rect 37001 42789 37013 42792
rect 37047 42789 37059 42823
rect 37001 42783 37059 42789
rect 27522 42752 27528 42764
rect 26988 42724 27528 42752
rect 26605 42715 26663 42721
rect 27522 42712 27528 42724
rect 27580 42712 27586 42764
rect 27893 42755 27951 42761
rect 27893 42721 27905 42755
rect 27939 42752 27951 42755
rect 28353 42755 28411 42761
rect 28353 42752 28365 42755
rect 27939 42724 28365 42752
rect 27939 42721 27951 42724
rect 27893 42715 27951 42721
rect 28353 42721 28365 42724
rect 28399 42721 28411 42755
rect 28353 42715 28411 42721
rect 28534 42712 28540 42764
rect 28592 42752 28598 42764
rect 30377 42755 30435 42761
rect 28592 42724 29776 42752
rect 28592 42712 28598 42724
rect 27249 42687 27307 42693
rect 27249 42684 27261 42687
rect 25740 42656 26188 42684
rect 26436 42656 27261 42684
rect 25740 42644 25746 42656
rect 26436 42548 26464 42656
rect 27249 42653 27261 42656
rect 27295 42684 27307 42687
rect 28074 42684 28080 42696
rect 27295 42656 28080 42684
rect 27295 42653 27307 42656
rect 27249 42647 27307 42653
rect 28074 42644 28080 42656
rect 28132 42644 28138 42696
rect 28442 42644 28448 42696
rect 28500 42684 28506 42696
rect 28905 42687 28963 42693
rect 28905 42684 28917 42687
rect 28500 42656 28917 42684
rect 28500 42644 28506 42656
rect 28905 42653 28917 42656
rect 28951 42653 28963 42687
rect 28905 42647 28963 42653
rect 29454 42644 29460 42696
rect 29512 42684 29518 42696
rect 29641 42687 29699 42693
rect 29641 42684 29653 42687
rect 29512 42656 29653 42684
rect 29512 42644 29518 42656
rect 29641 42653 29653 42656
rect 29687 42653 29699 42687
rect 29748 42684 29776 42724
rect 30377 42721 30389 42755
rect 30423 42752 30435 42755
rect 31018 42752 31024 42764
rect 30423 42724 31024 42752
rect 30423 42721 30435 42724
rect 30377 42715 30435 42721
rect 31018 42712 31024 42724
rect 31076 42712 31082 42764
rect 31294 42712 31300 42764
rect 31352 42752 31358 42764
rect 32217 42755 32275 42761
rect 31352 42724 32168 42752
rect 31352 42712 31358 42724
rect 30466 42684 30472 42696
rect 29748 42656 30472 42684
rect 29641 42647 29699 42653
rect 30466 42644 30472 42656
rect 30524 42644 30530 42696
rect 31665 42687 31723 42693
rect 31665 42653 31677 42687
rect 31711 42684 31723 42687
rect 31846 42684 31852 42696
rect 31711 42656 31852 42684
rect 31711 42653 31723 42656
rect 31665 42647 31723 42653
rect 31846 42644 31852 42656
rect 31904 42644 31910 42696
rect 32140 42684 32168 42724
rect 32217 42721 32229 42755
rect 32263 42752 32275 42755
rect 32306 42752 32312 42764
rect 32263 42724 32312 42752
rect 32263 42721 32275 42724
rect 32217 42715 32275 42721
rect 32306 42712 32312 42724
rect 32364 42712 32370 42764
rect 32508 42724 33456 42752
rect 32508 42693 32536 42724
rect 32493 42687 32551 42693
rect 32493 42684 32505 42687
rect 32140 42656 32505 42684
rect 32493 42653 32505 42656
rect 32539 42653 32551 42687
rect 32493 42647 32551 42653
rect 32585 42687 32643 42693
rect 32585 42653 32597 42687
rect 32631 42684 32643 42687
rect 33226 42684 33232 42696
rect 32631 42656 33232 42684
rect 32631 42653 32643 42656
rect 32585 42647 32643 42653
rect 33226 42644 33232 42656
rect 33284 42644 33290 42696
rect 33428 42628 33456 42724
rect 33502 42712 33508 42764
rect 33560 42712 33566 42764
rect 34054 42712 34060 42764
rect 34112 42752 34118 42764
rect 34425 42755 34483 42761
rect 34425 42752 34437 42755
rect 34112 42724 34437 42752
rect 34112 42712 34118 42724
rect 34425 42721 34437 42724
rect 34471 42721 34483 42755
rect 34425 42715 34483 42721
rect 36630 42712 36636 42764
rect 36688 42752 36694 42764
rect 37093 42755 37151 42761
rect 37093 42752 37105 42755
rect 36688 42724 37105 42752
rect 36688 42712 36694 42724
rect 37093 42721 37105 42724
rect 37139 42721 37151 42755
rect 37093 42715 37151 42721
rect 38102 42712 38108 42764
rect 38160 42752 38166 42764
rect 39577 42755 39635 42761
rect 38160 42724 39528 42752
rect 38160 42712 38166 42724
rect 33594 42644 33600 42696
rect 33652 42644 33658 42696
rect 33689 42687 33747 42693
rect 33689 42653 33701 42687
rect 33735 42653 33747 42687
rect 33689 42647 33747 42653
rect 34241 42687 34299 42693
rect 34241 42653 34253 42687
rect 34287 42684 34299 42687
rect 34974 42684 34980 42696
rect 34287 42656 34980 42684
rect 34287 42653 34299 42656
rect 34241 42647 34299 42653
rect 26510 42576 26516 42628
rect 26568 42616 26574 42628
rect 26568 42588 31754 42616
rect 26568 42576 26574 42588
rect 25056 42520 26464 42548
rect 24673 42511 24731 42517
rect 26694 42508 26700 42560
rect 26752 42508 26758 42560
rect 26878 42508 26884 42560
rect 26936 42548 26942 42560
rect 27525 42551 27583 42557
rect 27525 42548 27537 42551
rect 26936 42520 27537 42548
rect 26936 42508 26942 42520
rect 27525 42517 27537 42520
rect 27571 42517 27583 42551
rect 31726 42548 31754 42588
rect 32030 42576 32036 42628
rect 32088 42616 32094 42628
rect 33137 42619 33195 42625
rect 33137 42616 33149 42619
rect 32088 42588 33149 42616
rect 32088 42576 32094 42588
rect 33137 42585 33149 42588
rect 33183 42585 33195 42619
rect 33137 42579 33195 42585
rect 33410 42576 33416 42628
rect 33468 42616 33474 42628
rect 33704 42616 33732 42647
rect 34974 42644 34980 42656
rect 35032 42684 35038 42696
rect 35526 42684 35532 42696
rect 35032 42656 35532 42684
rect 35032 42644 35038 42656
rect 35526 42644 35532 42656
rect 35584 42684 35590 42696
rect 35897 42687 35955 42693
rect 35897 42684 35909 42687
rect 35584 42656 35909 42684
rect 35584 42644 35590 42656
rect 35897 42653 35909 42656
rect 35943 42653 35955 42687
rect 36814 42684 36820 42696
rect 35897 42647 35955 42653
rect 36004 42656 36820 42684
rect 33468 42588 33732 42616
rect 33468 42576 33474 42588
rect 35342 42576 35348 42628
rect 35400 42616 35406 42628
rect 36004 42616 36032 42656
rect 36814 42644 36820 42656
rect 36872 42644 36878 42696
rect 37182 42644 37188 42696
rect 37240 42684 37246 42696
rect 37553 42687 37611 42693
rect 37553 42684 37565 42687
rect 37240 42656 37565 42684
rect 37240 42644 37246 42656
rect 37553 42653 37565 42656
rect 37599 42653 37611 42687
rect 38378 42684 38384 42696
rect 37553 42647 37611 42653
rect 37660 42656 38384 42684
rect 35400 42588 36032 42616
rect 36541 42619 36599 42625
rect 35400 42576 35406 42588
rect 36541 42585 36553 42619
rect 36587 42616 36599 42619
rect 37660 42616 37688 42656
rect 38378 42644 38384 42656
rect 38436 42644 38442 42696
rect 38746 42644 38752 42696
rect 38804 42684 38810 42696
rect 38841 42687 38899 42693
rect 38841 42684 38853 42687
rect 38804 42656 38853 42684
rect 38804 42644 38810 42656
rect 38841 42653 38853 42656
rect 38887 42653 38899 42687
rect 39500 42684 39528 42724
rect 39577 42721 39589 42755
rect 39623 42752 39635 42755
rect 40144 42752 40172 42851
rect 40402 42848 40408 42900
rect 40460 42888 40466 42900
rect 40497 42891 40555 42897
rect 40497 42888 40509 42891
rect 40460 42860 40509 42888
rect 40460 42848 40466 42860
rect 40497 42857 40509 42860
rect 40543 42888 40555 42891
rect 41138 42888 41144 42900
rect 40543 42860 41144 42888
rect 40543 42857 40555 42860
rect 40497 42851 40555 42857
rect 41138 42848 41144 42860
rect 41196 42848 41202 42900
rect 41693 42891 41751 42897
rect 41693 42857 41705 42891
rect 41739 42888 41751 42891
rect 41966 42888 41972 42900
rect 41739 42860 41972 42888
rect 41739 42857 41751 42860
rect 41693 42851 41751 42857
rect 41966 42848 41972 42860
rect 42024 42848 42030 42900
rect 42518 42848 42524 42900
rect 42576 42848 42582 42900
rect 43990 42848 43996 42900
rect 44048 42888 44054 42900
rect 44085 42891 44143 42897
rect 44085 42888 44097 42891
rect 44048 42860 44097 42888
rect 44048 42848 44054 42860
rect 44085 42857 44097 42860
rect 44131 42857 44143 42891
rect 44085 42851 44143 42857
rect 46014 42848 46020 42900
rect 46072 42888 46078 42900
rect 46750 42888 46756 42900
rect 46072 42860 46756 42888
rect 46072 42848 46078 42860
rect 46750 42848 46756 42860
rect 46808 42848 46814 42900
rect 47394 42848 47400 42900
rect 47452 42888 47458 42900
rect 47857 42891 47915 42897
rect 47857 42888 47869 42891
rect 47452 42860 47869 42888
rect 47452 42848 47458 42860
rect 47857 42857 47869 42860
rect 47903 42857 47915 42891
rect 47857 42851 47915 42857
rect 48222 42848 48228 42900
rect 48280 42848 48286 42900
rect 51261 42891 51319 42897
rect 51261 42857 51273 42891
rect 51307 42888 51319 42891
rect 51534 42888 51540 42900
rect 51307 42860 51540 42888
rect 51307 42857 51319 42860
rect 51261 42851 51319 42857
rect 51534 42848 51540 42860
rect 51592 42848 51598 42900
rect 51629 42891 51687 42897
rect 51629 42857 51641 42891
rect 51675 42888 51687 42891
rect 52454 42888 52460 42900
rect 51675 42860 52460 42888
rect 51675 42857 51687 42860
rect 51629 42851 51687 42857
rect 52454 42848 52460 42860
rect 52512 42848 52518 42900
rect 41325 42823 41383 42829
rect 39623 42724 40172 42752
rect 40328 42792 41276 42820
rect 39623 42721 39635 42724
rect 39577 42715 39635 42721
rect 39669 42687 39727 42693
rect 39669 42684 39681 42687
rect 39500 42656 39681 42684
rect 38841 42647 38899 42653
rect 39669 42653 39681 42656
rect 39715 42684 39727 42687
rect 40328 42684 40356 42792
rect 39715 42656 40356 42684
rect 39715 42653 39727 42656
rect 39669 42647 39727 42653
rect 40586 42644 40592 42696
rect 40644 42644 40650 42696
rect 40770 42644 40776 42696
rect 40828 42644 40834 42696
rect 41064 42693 41092 42792
rect 41248 42752 41276 42792
rect 41325 42789 41337 42823
rect 41371 42820 41383 42823
rect 42536 42820 42564 42848
rect 41371 42792 42564 42820
rect 41371 42789 41383 42792
rect 41325 42783 41383 42789
rect 43162 42780 43168 42832
rect 43220 42780 43226 42832
rect 46658 42820 46664 42832
rect 46506 42792 46664 42820
rect 46658 42780 46664 42792
rect 46716 42780 46722 42832
rect 46842 42780 46848 42832
rect 46900 42780 46906 42832
rect 54018 42820 54024 42832
rect 53682 42792 54024 42820
rect 54018 42780 54024 42792
rect 54076 42780 54082 42832
rect 41414 42752 41420 42764
rect 41248 42724 41420 42752
rect 41414 42712 41420 42724
rect 41472 42752 41478 42764
rect 41782 42752 41788 42764
rect 41472 42724 41788 42752
rect 41472 42712 41478 42724
rect 41782 42712 41788 42724
rect 41840 42712 41846 42764
rect 44082 42712 44088 42764
rect 44140 42752 44146 42764
rect 46860 42752 46888 42780
rect 47305 42755 47363 42761
rect 47305 42752 47317 42755
rect 44140 42724 44312 42752
rect 46860 42724 47317 42752
rect 44140 42712 44146 42724
rect 41049 42687 41107 42693
rect 41049 42653 41061 42687
rect 41095 42653 41107 42687
rect 41049 42647 41107 42653
rect 41233 42687 41291 42693
rect 41233 42653 41245 42687
rect 41279 42684 41291 42687
rect 41279 42656 41736 42684
rect 41279 42653 41291 42656
rect 41233 42647 41291 42653
rect 36587 42588 37688 42616
rect 36587 42585 36599 42588
rect 36541 42579 36599 42585
rect 37826 42576 37832 42628
rect 37884 42616 37890 42628
rect 38289 42619 38347 42625
rect 38289 42616 38301 42619
rect 37884 42588 38301 42616
rect 37884 42576 37890 42588
rect 38289 42585 38301 42588
rect 38335 42585 38347 42619
rect 38289 42579 38347 42585
rect 38470 42576 38476 42628
rect 38528 42616 38534 42628
rect 41414 42616 41420 42628
rect 38528 42588 41420 42616
rect 38528 42576 38534 42588
rect 41414 42576 41420 42588
rect 41472 42576 41478 42628
rect 36446 42548 36452 42560
rect 31726 42520 36452 42548
rect 27525 42511 27583 42517
rect 36446 42508 36452 42520
rect 36504 42508 36510 42560
rect 37458 42508 37464 42560
rect 37516 42508 37522 42560
rect 38194 42508 38200 42560
rect 38252 42508 38258 42560
rect 38838 42508 38844 42560
rect 38896 42548 38902 42560
rect 39117 42551 39175 42557
rect 39117 42548 39129 42551
rect 38896 42520 39129 42548
rect 38896 42508 38902 42520
rect 39117 42517 39129 42520
rect 39163 42517 39175 42551
rect 39117 42511 39175 42517
rect 40034 42508 40040 42560
rect 40092 42548 40098 42560
rect 40586 42548 40592 42560
rect 40092 42520 40592 42548
rect 40092 42508 40098 42520
rect 40586 42508 40592 42520
rect 40644 42508 40650 42560
rect 41708 42548 41736 42656
rect 41874 42644 41880 42696
rect 41932 42644 41938 42696
rect 42150 42644 42156 42696
rect 42208 42644 42214 42696
rect 42518 42644 42524 42696
rect 42576 42684 42582 42696
rect 42576 42656 43760 42684
rect 42576 42644 42582 42656
rect 43732 42625 43760 42656
rect 44174 42644 44180 42696
rect 44232 42644 44238 42696
rect 44284 42693 44312 42724
rect 47305 42721 47317 42724
rect 47351 42721 47363 42755
rect 47305 42715 47363 42721
rect 47394 42712 47400 42764
rect 47452 42712 47458 42764
rect 48685 42755 48743 42761
rect 48685 42752 48697 42755
rect 47504 42724 48697 42752
rect 44269 42687 44327 42693
rect 44269 42653 44281 42687
rect 44315 42653 44327 42687
rect 44269 42647 44327 42653
rect 44910 42644 44916 42696
rect 44968 42684 44974 42696
rect 45005 42687 45063 42693
rect 45005 42684 45017 42687
rect 44968 42656 45017 42684
rect 44968 42644 44974 42656
rect 45005 42653 45017 42656
rect 45051 42653 45063 42687
rect 45005 42647 45063 42653
rect 45278 42644 45284 42696
rect 45336 42644 45342 42696
rect 46842 42644 46848 42696
rect 46900 42684 46906 42696
rect 47121 42687 47179 42693
rect 47121 42684 47133 42687
rect 46900 42656 47133 42684
rect 46900 42644 46906 42656
rect 47121 42653 47133 42656
rect 47167 42653 47179 42687
rect 47121 42647 47179 42653
rect 43717 42619 43775 42625
rect 43717 42585 43729 42619
rect 43763 42585 43775 42619
rect 43717 42579 43775 42585
rect 46290 42576 46296 42628
rect 46348 42616 46354 42628
rect 47504 42616 47532 42724
rect 48685 42721 48697 42724
rect 48731 42721 48743 42755
rect 48685 42715 48743 42721
rect 48317 42687 48375 42693
rect 48317 42684 48329 42687
rect 47780 42656 48329 42684
rect 47780 42625 47808 42656
rect 48317 42653 48329 42656
rect 48363 42653 48375 42687
rect 48317 42647 48375 42653
rect 48406 42644 48412 42696
rect 48464 42644 48470 42696
rect 49237 42687 49295 42693
rect 49237 42653 49249 42687
rect 49283 42653 49295 42687
rect 49237 42647 49295 42653
rect 46348 42588 47532 42616
rect 47765 42619 47823 42625
rect 46348 42576 46354 42588
rect 47765 42585 47777 42619
rect 47811 42585 47823 42619
rect 47765 42579 47823 42585
rect 43254 42548 43260 42560
rect 41708 42520 43260 42548
rect 43254 42508 43260 42520
rect 43312 42508 43318 42560
rect 43622 42508 43628 42560
rect 43680 42508 43686 42560
rect 46750 42508 46756 42560
rect 46808 42548 46814 42560
rect 49252 42548 49280 42647
rect 51718 42644 51724 42696
rect 51776 42644 51782 42696
rect 51902 42644 51908 42696
rect 51960 42644 51966 42696
rect 52181 42687 52239 42693
rect 52181 42653 52193 42687
rect 52227 42653 52239 42687
rect 52181 42647 52239 42653
rect 51534 42576 51540 42628
rect 51592 42616 51598 42628
rect 52196 42616 52224 42647
rect 52454 42644 52460 42696
rect 52512 42644 52518 42696
rect 52822 42644 52828 42696
rect 52880 42684 52886 42696
rect 54205 42687 54263 42693
rect 54205 42684 54217 42687
rect 52880 42656 54217 42684
rect 52880 42644 52886 42656
rect 54205 42653 54217 42656
rect 54251 42653 54263 42687
rect 54205 42647 54263 42653
rect 51592 42588 52224 42616
rect 51592 42576 51598 42588
rect 46808 42520 49280 42548
rect 46808 42508 46814 42520
rect 51902 42508 51908 42560
rect 51960 42548 51966 42560
rect 52914 42548 52920 42560
rect 51960 42520 52920 42548
rect 51960 42508 51966 42520
rect 52914 42508 52920 42520
rect 52972 42508 52978 42560
rect 552 42458 66424 42480
rect 552 42406 1998 42458
rect 2050 42406 2062 42458
rect 2114 42406 2126 42458
rect 2178 42406 2190 42458
rect 2242 42406 2254 42458
rect 2306 42406 49998 42458
rect 50050 42406 50062 42458
rect 50114 42406 50126 42458
rect 50178 42406 50190 42458
rect 50242 42406 50254 42458
rect 50306 42406 66424 42458
rect 552 42384 66424 42406
rect 11698 42304 11704 42356
rect 11756 42304 11762 42356
rect 12526 42304 12532 42356
rect 12584 42304 12590 42356
rect 15378 42304 15384 42356
rect 15436 42344 15442 42356
rect 16022 42344 16028 42356
rect 15436 42316 16028 42344
rect 15436 42304 15442 42316
rect 16022 42304 16028 42316
rect 16080 42304 16086 42356
rect 16298 42304 16304 42356
rect 16356 42344 16362 42356
rect 16356 42316 16712 42344
rect 16356 42304 16362 42316
rect 8386 42168 8392 42220
rect 8444 42208 8450 42220
rect 9953 42211 10011 42217
rect 9953 42208 9965 42211
rect 8444 42180 9965 42208
rect 8444 42168 8450 42180
rect 9953 42177 9965 42180
rect 9999 42208 10011 42211
rect 11514 42208 11520 42220
rect 9999 42180 11520 42208
rect 9999 42177 10011 42180
rect 9953 42171 10011 42177
rect 11514 42168 11520 42180
rect 11572 42168 11578 42220
rect 12986 42168 12992 42220
rect 13044 42168 13050 42220
rect 13170 42168 13176 42220
rect 13228 42168 13234 42220
rect 15396 42217 15424 42304
rect 16684 42276 16712 42316
rect 16942 42304 16948 42356
rect 17000 42344 17006 42356
rect 17589 42347 17647 42353
rect 17589 42344 17601 42347
rect 17000 42316 17601 42344
rect 17000 42304 17006 42316
rect 17589 42313 17601 42316
rect 17635 42313 17647 42347
rect 17589 42307 17647 42313
rect 17862 42304 17868 42356
rect 17920 42344 17926 42356
rect 17920 42316 18184 42344
rect 17920 42304 17926 42316
rect 17954 42276 17960 42288
rect 16684 42248 17960 42276
rect 17954 42236 17960 42248
rect 18012 42236 18018 42288
rect 15381 42211 15439 42217
rect 15381 42177 15393 42211
rect 15427 42177 15439 42211
rect 15381 42171 15439 42177
rect 15657 42211 15715 42217
rect 15657 42177 15669 42211
rect 15703 42208 15715 42211
rect 16390 42208 16396 42220
rect 15703 42180 16396 42208
rect 15703 42177 15715 42180
rect 15657 42171 15715 42177
rect 16390 42168 16396 42180
rect 16448 42168 16454 42220
rect 16666 42168 16672 42220
rect 16724 42208 16730 42220
rect 16724 42180 17816 42208
rect 16724 42168 16730 42180
rect 9674 42100 9680 42152
rect 9732 42100 9738 42152
rect 13722 42100 13728 42152
rect 13780 42100 13786 42152
rect 14553 42143 14611 42149
rect 14553 42109 14565 42143
rect 14599 42109 14611 42143
rect 17678 42140 17684 42152
rect 16790 42112 17684 42140
rect 14553 42103 14611 42109
rect 10229 42075 10287 42081
rect 10229 42041 10241 42075
rect 10275 42041 10287 42075
rect 11977 42075 12035 42081
rect 11977 42072 11989 42075
rect 11454 42044 11989 42072
rect 10229 42035 10287 42041
rect 11977 42041 11989 42044
rect 12023 42041 12035 42075
rect 11977 42035 12035 42041
rect 8570 41964 8576 42016
rect 8628 42004 8634 42016
rect 9033 42007 9091 42013
rect 9033 42004 9045 42007
rect 8628 41976 9045 42004
rect 8628 41964 8634 41976
rect 9033 41973 9045 41976
rect 9079 41973 9091 42007
rect 10244 42004 10272 42035
rect 11054 42004 11060 42016
rect 10244 41976 11060 42004
rect 9033 41967 9091 41973
rect 11054 41964 11060 41976
rect 11112 41964 11118 42016
rect 11992 42004 12020 42035
rect 12250 42032 12256 42084
rect 12308 42072 12314 42084
rect 12345 42075 12403 42081
rect 12345 42072 12357 42075
rect 12308 42044 12357 42072
rect 12308 42032 12314 42044
rect 12345 42041 12357 42044
rect 12391 42041 12403 42075
rect 12345 42035 12403 42041
rect 12710 42032 12716 42084
rect 12768 42072 12774 42084
rect 12897 42075 12955 42081
rect 12897 42072 12909 42075
rect 12768 42044 12909 42072
rect 12768 42032 12774 42044
rect 12897 42041 12909 42044
rect 12943 42072 12955 42075
rect 13630 42072 13636 42084
rect 12943 42044 13636 42072
rect 12943 42041 12955 42044
rect 12897 42035 12955 42041
rect 13630 42032 13636 42044
rect 13688 42032 13694 42084
rect 14568 42072 14596 42103
rect 17678 42100 17684 42112
rect 17736 42100 17742 42152
rect 17788 42140 17816 42180
rect 18046 42168 18052 42220
rect 18104 42168 18110 42220
rect 18156 42217 18184 42316
rect 19794 42304 19800 42356
rect 19852 42304 19858 42356
rect 20165 42347 20223 42353
rect 20165 42313 20177 42347
rect 20211 42344 20223 42347
rect 20438 42344 20444 42356
rect 20211 42316 20444 42344
rect 20211 42313 20223 42316
rect 20165 42307 20223 42313
rect 20438 42304 20444 42316
rect 20496 42304 20502 42356
rect 24762 42304 24768 42356
rect 24820 42304 24826 42356
rect 24946 42304 24952 42356
rect 25004 42344 25010 42356
rect 25593 42347 25651 42353
rect 25004 42316 25360 42344
rect 25004 42304 25010 42316
rect 22097 42279 22155 42285
rect 22097 42245 22109 42279
rect 22143 42276 22155 42279
rect 22278 42276 22284 42288
rect 22143 42248 22284 42276
rect 22143 42245 22155 42248
rect 22097 42239 22155 42245
rect 22278 42236 22284 42248
rect 22336 42236 22342 42288
rect 25222 42276 25228 42288
rect 23584 42248 25228 42276
rect 18141 42211 18199 42217
rect 18141 42177 18153 42211
rect 18187 42208 18199 42211
rect 19153 42211 19211 42217
rect 19153 42208 19165 42211
rect 18187 42180 19165 42208
rect 18187 42177 18199 42180
rect 18141 42171 18199 42177
rect 19153 42177 19165 42180
rect 19199 42208 19211 42211
rect 20530 42208 20536 42220
rect 19199 42180 20536 42208
rect 19199 42177 19211 42180
rect 19153 42171 19211 42177
rect 20530 42168 20536 42180
rect 20588 42168 20594 42220
rect 22002 42168 22008 42220
rect 22060 42168 22066 42220
rect 22554 42168 22560 42220
rect 22612 42168 22618 42220
rect 23584 42217 23612 42248
rect 25222 42236 25228 42248
rect 25280 42236 25286 42288
rect 25332 42276 25360 42316
rect 25593 42313 25605 42347
rect 25639 42344 25651 42347
rect 25958 42344 25964 42356
rect 25639 42316 25964 42344
rect 25639 42313 25651 42316
rect 25593 42307 25651 42313
rect 25958 42304 25964 42316
rect 26016 42304 26022 42356
rect 28350 42304 28356 42356
rect 28408 42304 28414 42356
rect 32879 42347 32937 42353
rect 32879 42313 32891 42347
rect 32925 42344 32937 42347
rect 33042 42344 33048 42356
rect 32925 42316 33048 42344
rect 32925 42313 32937 42316
rect 32879 42307 32937 42313
rect 33042 42304 33048 42316
rect 33100 42304 33106 42356
rect 33226 42304 33232 42356
rect 33284 42304 33290 42356
rect 33502 42304 33508 42356
rect 33560 42344 33566 42356
rect 34149 42347 34207 42353
rect 34149 42344 34161 42347
rect 33560 42316 34161 42344
rect 33560 42304 33566 42316
rect 34149 42313 34161 42316
rect 34195 42313 34207 42347
rect 34149 42307 34207 42313
rect 35897 42347 35955 42353
rect 35897 42313 35909 42347
rect 35943 42344 35955 42347
rect 36170 42344 36176 42356
rect 35943 42316 36176 42344
rect 35943 42313 35955 42316
rect 35897 42307 35955 42313
rect 36170 42304 36176 42316
rect 36228 42304 36234 42356
rect 36446 42304 36452 42356
rect 36504 42344 36510 42356
rect 36504 42316 40632 42344
rect 36504 42304 36510 42316
rect 25332 42248 26280 42276
rect 22649 42211 22707 42217
rect 22649 42177 22661 42211
rect 22695 42177 22707 42211
rect 22649 42171 22707 42177
rect 23569 42211 23627 42217
rect 23569 42177 23581 42211
rect 23615 42177 23627 42211
rect 23569 42171 23627 42177
rect 18322 42140 18328 42152
rect 17788 42112 18328 42140
rect 18322 42100 18328 42112
rect 18380 42100 18386 42152
rect 19334 42100 19340 42152
rect 19392 42140 19398 42152
rect 19429 42143 19487 42149
rect 19429 42140 19441 42143
rect 19392 42112 19441 42140
rect 19392 42100 19398 42112
rect 19429 42109 19441 42112
rect 19475 42109 19487 42143
rect 19429 42103 19487 42109
rect 22094 42100 22100 42152
rect 22152 42140 22158 42152
rect 22465 42143 22523 42149
rect 22465 42140 22477 42143
rect 22152 42112 22477 42140
rect 22152 42100 22158 42112
rect 22465 42109 22477 42112
rect 22511 42109 22523 42143
rect 22465 42103 22523 42109
rect 17497 42075 17555 42081
rect 14568 42044 16068 42072
rect 12434 42004 12440 42016
rect 11992 41976 12440 42004
rect 12434 41964 12440 41976
rect 12492 41964 12498 42016
rect 14366 41964 14372 42016
rect 14424 41964 14430 42016
rect 15105 42007 15163 42013
rect 15105 41973 15117 42007
rect 15151 42004 15163 42007
rect 15470 42004 15476 42016
rect 15151 41976 15476 42004
rect 15151 41973 15163 41976
rect 15105 41967 15163 41973
rect 15470 41964 15476 41976
rect 15528 41964 15534 42016
rect 16040 42004 16068 42044
rect 17497 42041 17509 42075
rect 17543 42072 17555 42075
rect 17954 42072 17960 42084
rect 17543 42044 17960 42072
rect 17543 42041 17555 42044
rect 17497 42035 17555 42041
rect 17954 42032 17960 42044
rect 18012 42032 18018 42084
rect 20438 42032 20444 42084
rect 20496 42072 20502 42084
rect 20496 42044 20562 42072
rect 20496 42032 20502 42044
rect 21450 42032 21456 42084
rect 21508 42072 21514 42084
rect 21729 42075 21787 42081
rect 21729 42072 21741 42075
rect 21508 42044 21741 42072
rect 21508 42032 21514 42044
rect 21729 42041 21741 42044
rect 21775 42041 21787 42075
rect 21729 42035 21787 42041
rect 21818 42032 21824 42084
rect 21876 42072 21882 42084
rect 22664 42072 22692 42171
rect 24026 42168 24032 42220
rect 24084 42208 24090 42220
rect 26252 42217 26280 42248
rect 28074 42236 28080 42288
rect 28132 42276 28138 42288
rect 28810 42276 28816 42288
rect 28132 42248 28816 42276
rect 28132 42236 28138 42248
rect 28810 42236 28816 42248
rect 28868 42236 28874 42288
rect 35342 42276 35348 42288
rect 33796 42248 35348 42276
rect 24121 42211 24179 42217
rect 24121 42208 24133 42211
rect 24084 42180 24133 42208
rect 24084 42168 24090 42180
rect 24121 42177 24133 42180
rect 24167 42177 24179 42211
rect 26145 42211 26203 42217
rect 26145 42208 26157 42211
rect 24121 42171 24179 42177
rect 24228 42180 26157 42208
rect 23014 42100 23020 42152
rect 23072 42140 23078 42152
rect 23293 42143 23351 42149
rect 23293 42140 23305 42143
rect 23072 42112 23305 42140
rect 23072 42100 23078 42112
rect 23293 42109 23305 42112
rect 23339 42109 23351 42143
rect 23293 42103 23351 42109
rect 23385 42143 23443 42149
rect 23385 42109 23397 42143
rect 23431 42140 23443 42143
rect 23431 42112 23704 42140
rect 23431 42109 23443 42112
rect 23385 42103 23443 42109
rect 21876 42044 22692 42072
rect 23676 42072 23704 42112
rect 23750 42100 23756 42152
rect 23808 42140 23814 42152
rect 24228 42140 24256 42180
rect 26145 42177 26157 42180
rect 26191 42177 26203 42211
rect 26145 42171 26203 42177
rect 26237 42211 26295 42217
rect 26237 42177 26249 42211
rect 26283 42177 26295 42211
rect 26237 42171 26295 42177
rect 26602 42168 26608 42220
rect 26660 42168 26666 42220
rect 27430 42168 27436 42220
rect 27488 42208 27494 42220
rect 32122 42208 32128 42220
rect 27488 42180 32128 42208
rect 27488 42168 27494 42180
rect 32122 42168 32128 42180
rect 32180 42168 32186 42220
rect 32214 42168 32220 42220
rect 32272 42208 32278 42220
rect 33137 42211 33195 42217
rect 33137 42208 33149 42211
rect 32272 42180 33149 42208
rect 32272 42168 32278 42180
rect 33137 42177 33149 42180
rect 33183 42177 33195 42211
rect 33137 42171 33195 42177
rect 33226 42168 33232 42220
rect 33284 42208 33290 42220
rect 33796 42217 33824 42248
rect 35342 42236 35348 42248
rect 35400 42236 35406 42288
rect 33781 42211 33839 42217
rect 33781 42208 33793 42211
rect 33284 42180 33793 42208
rect 33284 42168 33290 42180
rect 33781 42177 33793 42180
rect 33827 42177 33839 42211
rect 33781 42171 33839 42177
rect 34422 42168 34428 42220
rect 34480 42208 34486 42220
rect 34701 42211 34759 42217
rect 34701 42208 34713 42211
rect 34480 42180 34713 42208
rect 34480 42168 34486 42180
rect 34701 42177 34713 42180
rect 34747 42177 34759 42211
rect 34701 42171 34759 42177
rect 37458 42168 37464 42220
rect 37516 42208 37522 42220
rect 38289 42211 38347 42217
rect 38289 42208 38301 42211
rect 37516 42180 38301 42208
rect 37516 42168 37522 42180
rect 38289 42177 38301 42180
rect 38335 42177 38347 42211
rect 38289 42171 38347 42177
rect 38378 42168 38384 42220
rect 38436 42168 38442 42220
rect 39301 42211 39359 42217
rect 39301 42177 39313 42211
rect 39347 42208 39359 42211
rect 40310 42208 40316 42220
rect 39347 42180 40316 42208
rect 39347 42177 39359 42180
rect 39301 42171 39359 42177
rect 40310 42168 40316 42180
rect 40368 42168 40374 42220
rect 40604 42208 40632 42316
rect 40770 42304 40776 42356
rect 40828 42344 40834 42356
rect 41233 42347 41291 42353
rect 41233 42344 41245 42347
rect 40828 42316 41245 42344
rect 40828 42304 40834 42316
rect 41233 42313 41245 42316
rect 41279 42344 41291 42347
rect 43898 42344 43904 42356
rect 41279 42316 43904 42344
rect 41279 42313 41291 42316
rect 41233 42307 41291 42313
rect 43898 42304 43904 42316
rect 43956 42304 43962 42356
rect 44266 42304 44272 42356
rect 44324 42344 44330 42356
rect 44453 42347 44511 42353
rect 44453 42344 44465 42347
rect 44324 42316 44465 42344
rect 44324 42304 44330 42316
rect 44453 42313 44465 42316
rect 44499 42313 44511 42347
rect 44453 42307 44511 42313
rect 45278 42304 45284 42356
rect 45336 42344 45342 42356
rect 45557 42347 45615 42353
rect 45557 42344 45569 42347
rect 45336 42316 45569 42344
rect 45336 42304 45342 42316
rect 45557 42313 45569 42316
rect 45603 42313 45615 42347
rect 45557 42307 45615 42313
rect 49694 42304 49700 42356
rect 49752 42344 49758 42356
rect 51626 42344 51632 42356
rect 49752 42316 51632 42344
rect 49752 42304 49758 42316
rect 45922 42276 45928 42288
rect 41386 42248 45928 42276
rect 41386 42208 41414 42248
rect 45922 42236 45928 42248
rect 45980 42236 45986 42288
rect 40604 42180 41414 42208
rect 44082 42168 44088 42220
rect 44140 42208 44146 42220
rect 45005 42211 45063 42217
rect 45005 42208 45017 42211
rect 44140 42180 45017 42208
rect 44140 42168 44146 42180
rect 45005 42177 45017 42180
rect 45051 42177 45063 42211
rect 45005 42171 45063 42177
rect 45830 42168 45836 42220
rect 45888 42208 45894 42220
rect 46109 42211 46167 42217
rect 46109 42208 46121 42211
rect 45888 42180 46121 42208
rect 45888 42168 45894 42180
rect 46109 42177 46121 42180
rect 46155 42208 46167 42211
rect 46750 42208 46756 42220
rect 46155 42180 46756 42208
rect 46155 42177 46167 42180
rect 46109 42171 46167 42177
rect 46750 42168 46756 42180
rect 46808 42168 46814 42220
rect 47762 42168 47768 42220
rect 47820 42208 47826 42220
rect 48225 42211 48283 42217
rect 48225 42208 48237 42211
rect 47820 42180 48237 42208
rect 47820 42168 47826 42180
rect 48225 42177 48237 42180
rect 48271 42208 48283 42211
rect 48409 42211 48467 42217
rect 48409 42208 48421 42211
rect 48271 42180 48421 42208
rect 48271 42177 48283 42180
rect 48225 42171 48283 42177
rect 48409 42177 48421 42180
rect 48455 42177 48467 42211
rect 48409 42171 48467 42177
rect 49142 42168 49148 42220
rect 49200 42208 49206 42220
rect 51000 42217 51028 42316
rect 51626 42304 51632 42316
rect 51684 42304 51690 42356
rect 51718 42304 51724 42356
rect 51776 42344 51782 42356
rect 51997 42347 52055 42353
rect 51997 42344 52009 42347
rect 51776 42316 52009 42344
rect 51776 42304 51782 42316
rect 51997 42313 52009 42316
rect 52043 42313 52055 42347
rect 51997 42307 52055 42313
rect 52089 42347 52147 42353
rect 52089 42313 52101 42347
rect 52135 42344 52147 42347
rect 52454 42344 52460 42356
rect 52135 42316 52460 42344
rect 52135 42313 52147 42316
rect 52089 42307 52147 42313
rect 52454 42304 52460 42316
rect 52512 42304 52518 42356
rect 53190 42304 53196 42356
rect 53248 42344 53254 42356
rect 59262 42344 59268 42356
rect 53248 42316 59268 42344
rect 53248 42304 53254 42316
rect 59262 42304 59268 42316
rect 59320 42304 59326 42356
rect 53101 42279 53159 42285
rect 53101 42276 53113 42279
rect 51644 42248 53113 42276
rect 50157 42211 50215 42217
rect 50157 42208 50169 42211
rect 49200 42180 50169 42208
rect 49200 42168 49206 42180
rect 50157 42177 50169 42180
rect 50203 42177 50215 42211
rect 50157 42171 50215 42177
rect 50985 42211 51043 42217
rect 50985 42177 50997 42211
rect 51031 42177 51043 42211
rect 50985 42171 51043 42177
rect 51445 42211 51503 42217
rect 51445 42177 51457 42211
rect 51491 42208 51503 42211
rect 51644 42208 51672 42248
rect 53101 42245 53113 42248
rect 53147 42276 53159 42279
rect 53147 42248 53328 42276
rect 53147 42245 53159 42248
rect 53101 42239 53159 42245
rect 51491 42180 51672 42208
rect 51491 42177 51503 42180
rect 51445 42171 51503 42177
rect 51718 42168 51724 42220
rect 51776 42208 51782 42220
rect 52638 42208 52644 42220
rect 51776 42180 52644 42208
rect 51776 42168 51782 42180
rect 52638 42168 52644 42180
rect 52696 42168 52702 42220
rect 53300 42208 53328 42248
rect 53374 42236 53380 42288
rect 53432 42276 53438 42288
rect 62666 42276 62672 42288
rect 53432 42248 62672 42276
rect 53432 42236 53438 42248
rect 62666 42236 62672 42248
rect 62724 42236 62730 42288
rect 53926 42208 53932 42220
rect 53300 42180 53932 42208
rect 53926 42168 53932 42180
rect 53984 42168 53990 42220
rect 23808 42112 24256 42140
rect 24305 42143 24363 42149
rect 23808 42100 23814 42112
rect 24305 42109 24317 42143
rect 24351 42140 24363 42143
rect 25038 42140 25044 42152
rect 24351 42112 25044 42140
rect 24351 42109 24363 42112
rect 24305 42103 24363 42109
rect 25038 42100 25044 42112
rect 25096 42140 25102 42152
rect 26053 42143 26111 42149
rect 26053 42140 26065 42143
rect 25096 42112 26065 42140
rect 25096 42100 25102 42112
rect 26053 42109 26065 42112
rect 26099 42109 26111 42143
rect 28442 42140 28448 42152
rect 28014 42112 28448 42140
rect 26053 42103 26111 42109
rect 28442 42100 28448 42112
rect 28500 42140 28506 42152
rect 29086 42140 29092 42152
rect 28500 42112 29092 42140
rect 28500 42100 28506 42112
rect 29086 42100 29092 42112
rect 29144 42140 29150 42152
rect 29365 42143 29423 42149
rect 29365 42140 29377 42143
rect 29144 42112 29377 42140
rect 29144 42100 29150 42112
rect 29365 42109 29377 42112
rect 29411 42109 29423 42143
rect 29365 42103 29423 42109
rect 31754 42100 31760 42152
rect 31812 42100 31818 42152
rect 33597 42143 33655 42149
rect 33597 42109 33609 42143
rect 33643 42140 33655 42143
rect 34440 42140 34468 42168
rect 33643 42112 34468 42140
rect 33643 42109 33655 42112
rect 33597 42103 33655 42109
rect 35066 42100 35072 42152
rect 35124 42140 35130 42152
rect 35618 42140 35624 42152
rect 35124 42112 35624 42140
rect 35124 42100 35130 42112
rect 35618 42100 35624 42112
rect 35676 42100 35682 42152
rect 37734 42100 37740 42152
rect 37792 42100 37798 42152
rect 38194 42100 38200 42152
rect 38252 42100 38258 42152
rect 41414 42100 41420 42152
rect 41472 42140 41478 42152
rect 41472 42112 41920 42140
rect 41472 42100 41478 42112
rect 41892 42084 41920 42112
rect 44450 42100 44456 42152
rect 44508 42140 44514 42152
rect 44913 42143 44971 42149
rect 44913 42140 44925 42143
rect 44508 42112 44925 42140
rect 44508 42100 44514 42112
rect 44913 42109 44925 42112
rect 44959 42109 44971 42143
rect 44913 42103 44971 42109
rect 45094 42100 45100 42152
rect 45152 42140 45158 42152
rect 46477 42143 46535 42149
rect 46477 42140 46489 42143
rect 45152 42112 46489 42140
rect 45152 42100 45158 42112
rect 46477 42109 46489 42112
rect 46523 42109 46535 42143
rect 46477 42103 46535 42109
rect 49973 42143 50031 42149
rect 49973 42109 49985 42143
rect 50019 42140 50031 42143
rect 52362 42140 52368 42152
rect 50019 42112 52368 42140
rect 50019 42109 50031 42112
rect 49973 42103 50031 42109
rect 52362 42100 52368 42112
rect 52420 42100 52426 42152
rect 52457 42143 52515 42149
rect 52457 42109 52469 42143
rect 52503 42140 52515 42143
rect 52546 42140 52552 42152
rect 52503 42112 52552 42140
rect 52503 42109 52515 42112
rect 52457 42103 52515 42109
rect 52546 42100 52552 42112
rect 52604 42100 52610 42152
rect 53374 42100 53380 42152
rect 53432 42100 53438 42152
rect 53834 42100 53840 42152
rect 53892 42140 53898 42152
rect 63034 42140 63040 42152
rect 53892 42112 63040 42140
rect 53892 42100 53898 42112
rect 63034 42100 63040 42112
rect 63092 42100 63098 42152
rect 23676 42044 25728 42072
rect 21876 42032 21882 42044
rect 17034 42004 17040 42016
rect 16040 41976 17040 42004
rect 17034 41964 17040 41976
rect 17092 41964 17098 42016
rect 17129 42007 17187 42013
rect 17129 41973 17141 42007
rect 17175 42004 17187 42007
rect 17218 42004 17224 42016
rect 17175 41976 17224 42004
rect 17175 41973 17187 41976
rect 17129 41967 17187 41973
rect 17218 41964 17224 41976
rect 17276 41964 17282 42016
rect 17586 41964 17592 42016
rect 17644 42004 17650 42016
rect 17862 42004 17868 42016
rect 17644 41976 17868 42004
rect 17644 41964 17650 41976
rect 17862 41964 17868 41976
rect 17920 41964 17926 42016
rect 19337 42007 19395 42013
rect 19337 41973 19349 42007
rect 19383 42004 19395 42007
rect 19702 42004 19708 42016
rect 19383 41976 19708 42004
rect 19383 41973 19395 41976
rect 19337 41967 19395 41973
rect 19702 41964 19708 41976
rect 19760 41964 19766 42016
rect 20257 42007 20315 42013
rect 20257 41973 20269 42007
rect 20303 42004 20315 42007
rect 22278 42004 22284 42016
rect 20303 41976 22284 42004
rect 20303 41973 20315 41976
rect 20257 41967 20315 41973
rect 22278 41964 22284 41976
rect 22336 42004 22342 42016
rect 22738 42004 22744 42016
rect 22336 41976 22744 42004
rect 22336 41964 22342 41976
rect 22738 41964 22744 41976
rect 22796 41964 22802 42016
rect 22925 42007 22983 42013
rect 22925 41973 22937 42007
rect 22971 42004 22983 42007
rect 23290 42004 23296 42016
rect 22971 41976 23296 42004
rect 22971 41973 22983 41976
rect 22925 41967 22983 41973
rect 23290 41964 23296 41976
rect 23348 41964 23354 42016
rect 24397 42007 24455 42013
rect 24397 41973 24409 42007
rect 24443 42004 24455 42007
rect 25406 42004 25412 42016
rect 24443 41976 25412 42004
rect 24443 41973 24455 41976
rect 24397 41967 24455 41973
rect 25406 41964 25412 41976
rect 25464 41964 25470 42016
rect 25700 42013 25728 42044
rect 26878 42032 26884 42084
rect 26936 42032 26942 42084
rect 28184 42044 29224 42072
rect 25685 42007 25743 42013
rect 25685 41973 25697 42007
rect 25731 41973 25743 42007
rect 25685 41967 25743 41973
rect 25774 41964 25780 42016
rect 25832 42004 25838 42016
rect 28184 42004 28212 42044
rect 25832 41976 28212 42004
rect 25832 41964 25838 41976
rect 28258 41964 28264 42016
rect 28316 42004 28322 42016
rect 29089 42007 29147 42013
rect 29089 42004 29101 42007
rect 28316 41976 29101 42004
rect 28316 41964 28322 41976
rect 29089 41973 29101 41976
rect 29135 41973 29147 42007
rect 29196 42004 29224 42044
rect 32858 42032 32864 42084
rect 32916 42072 32922 42084
rect 35894 42072 35900 42084
rect 32916 42044 35900 42072
rect 32916 42032 32922 42044
rect 35894 42032 35900 42044
rect 35952 42032 35958 42084
rect 36078 42032 36084 42084
rect 36136 42072 36142 42084
rect 37461 42075 37519 42081
rect 36136 42044 36294 42072
rect 36136 42032 36142 42044
rect 37461 42041 37473 42075
rect 37507 42072 37519 42075
rect 37507 42044 37872 42072
rect 37507 42041 37519 42044
rect 37461 42035 37519 42041
rect 30374 42004 30380 42016
rect 29196 41976 30380 42004
rect 29089 41967 29147 41973
rect 30374 41964 30380 41976
rect 30432 41964 30438 42016
rect 31389 42007 31447 42013
rect 31389 41973 31401 42007
rect 31435 42004 31447 42007
rect 31846 42004 31852 42016
rect 31435 41976 31852 42004
rect 31435 41973 31447 41976
rect 31389 41967 31447 41973
rect 31846 41964 31852 41976
rect 31904 42004 31910 42016
rect 33226 42004 33232 42016
rect 31904 41976 33232 42004
rect 31904 41964 31910 41976
rect 33226 41964 33232 41976
rect 33284 41964 33290 42016
rect 33689 42007 33747 42013
rect 33689 41973 33701 42007
rect 33735 42004 33747 42007
rect 33778 42004 33784 42016
rect 33735 41976 33784 42004
rect 33735 41973 33747 41976
rect 33689 41967 33747 41973
rect 33778 41964 33784 41976
rect 33836 41964 33842 42016
rect 35989 42007 36047 42013
rect 35989 41973 36001 42007
rect 36035 42004 36047 42007
rect 37182 42004 37188 42016
rect 36035 41976 37188 42004
rect 36035 41973 36047 41976
rect 35989 41967 36047 41973
rect 37182 41964 37188 41976
rect 37240 41964 37246 42016
rect 37844 42013 37872 42044
rect 39574 42032 39580 42084
rect 39632 42032 39638 42084
rect 40954 42072 40960 42084
rect 40802 42044 40960 42072
rect 40954 42032 40960 42044
rect 41012 42032 41018 42084
rect 41506 42032 41512 42084
rect 41564 42032 41570 42084
rect 41874 42032 41880 42084
rect 41932 42032 41938 42084
rect 43162 42032 43168 42084
rect 43220 42072 43226 42084
rect 43220 42044 43392 42072
rect 43220 42032 43226 42044
rect 37829 42007 37887 42013
rect 37829 41973 37841 42007
rect 37875 41973 37887 42007
rect 37829 41967 37887 41973
rect 41049 42007 41107 42013
rect 41049 41973 41061 42007
rect 41095 42004 41107 42007
rect 41138 42004 41144 42016
rect 41095 41976 41144 42004
rect 41095 41973 41107 41976
rect 41049 41967 41107 41973
rect 41138 41964 41144 41976
rect 41196 41964 41202 42016
rect 43364 42004 43392 42044
rect 43438 42032 43444 42084
rect 43496 42072 43502 42084
rect 43625 42075 43683 42081
rect 43625 42072 43637 42075
rect 43496 42044 43637 42072
rect 43496 42032 43502 42044
rect 43625 42041 43637 42044
rect 43671 42041 43683 42075
rect 43625 42035 43683 42041
rect 44266 42032 44272 42084
rect 44324 42072 44330 42084
rect 44821 42075 44879 42081
rect 44821 42072 44833 42075
rect 44324 42044 44833 42072
rect 44324 42032 44330 42044
rect 44821 42041 44833 42044
rect 44867 42072 44879 42075
rect 45281 42075 45339 42081
rect 45281 42072 45293 42075
rect 44867 42044 45293 42072
rect 44867 42041 44879 42044
rect 44821 42035 44879 42041
rect 45281 42041 45293 42044
rect 45327 42041 45339 42075
rect 45281 42035 45339 42041
rect 45925 42075 45983 42081
rect 45925 42041 45937 42075
rect 45971 42072 45983 42075
rect 46290 42072 46296 42084
rect 45971 42044 46296 42072
rect 45971 42041 45983 42044
rect 45925 42035 45983 42041
rect 46290 42032 46296 42044
rect 46348 42032 46354 42084
rect 46753 42075 46811 42081
rect 46753 42041 46765 42075
rect 46799 42041 46811 42075
rect 48038 42072 48044 42084
rect 47978 42044 48044 42072
rect 46753 42035 46811 42041
rect 45830 42004 45836 42016
rect 43364 41976 45836 42004
rect 45830 41964 45836 41976
rect 45888 41964 45894 42016
rect 46014 41964 46020 42016
rect 46072 41964 46078 42016
rect 46768 42004 46796 42035
rect 48038 42032 48044 42044
rect 48096 42072 48102 42084
rect 48314 42072 48320 42084
rect 48096 42044 48320 42072
rect 48096 42032 48102 42044
rect 48314 42032 48320 42044
rect 48372 42032 48378 42084
rect 49878 42032 49884 42084
rect 49936 42072 49942 42084
rect 50065 42075 50123 42081
rect 50065 42072 50077 42075
rect 49936 42044 50077 42072
rect 49936 42032 49942 42044
rect 50065 42041 50077 42044
rect 50111 42041 50123 42075
rect 50065 42035 50123 42041
rect 50801 42075 50859 42081
rect 50801 42041 50813 42075
rect 50847 42072 50859 42075
rect 51350 42072 51356 42084
rect 50847 42044 51356 42072
rect 50847 42041 50859 42044
rect 50801 42035 50859 42041
rect 51350 42032 51356 42044
rect 51408 42032 51414 42084
rect 53190 42032 53196 42084
rect 53248 42072 53254 42084
rect 53653 42075 53711 42081
rect 53653 42072 53665 42075
rect 53248 42044 53665 42072
rect 53248 42032 53254 42044
rect 53653 42041 53665 42044
rect 53699 42041 53711 42075
rect 53653 42035 53711 42041
rect 54018 42032 54024 42084
rect 54076 42032 54082 42084
rect 55766 42032 55772 42084
rect 55824 42032 55830 42084
rect 48130 42004 48136 42016
rect 46768 41976 48136 42004
rect 48130 41964 48136 41976
rect 48188 41964 48194 42016
rect 48498 41964 48504 42016
rect 48556 42004 48562 42016
rect 49053 42007 49111 42013
rect 49053 42004 49065 42007
rect 48556 41976 49065 42004
rect 48556 41964 48562 41976
rect 49053 41973 49065 41976
rect 49099 41973 49111 42007
rect 49053 41967 49111 41973
rect 49605 42007 49663 42013
rect 49605 41973 49617 42007
rect 49651 42004 49663 42007
rect 49786 42004 49792 42016
rect 49651 41976 49792 42004
rect 49651 41973 49663 41976
rect 49605 41967 49663 41973
rect 49786 41964 49792 41976
rect 49844 41964 49850 42016
rect 50430 41964 50436 42016
rect 50488 41964 50494 42016
rect 50706 41964 50712 42016
rect 50764 42004 50770 42016
rect 50893 42007 50951 42013
rect 50893 42004 50905 42007
rect 50764 41976 50905 42004
rect 50764 41964 50770 41976
rect 50893 41973 50905 41976
rect 50939 42004 50951 42007
rect 51537 42007 51595 42013
rect 51537 42004 51549 42007
rect 50939 41976 51549 42004
rect 50939 41973 50951 41976
rect 50893 41967 50951 41973
rect 51537 41973 51549 41976
rect 51583 41973 51595 42007
rect 51537 41967 51595 41973
rect 51629 42007 51687 42013
rect 51629 41973 51641 42007
rect 51675 42004 51687 42007
rect 52454 42004 52460 42016
rect 51675 41976 52460 42004
rect 51675 41973 51687 41976
rect 51629 41967 51687 41973
rect 52454 41964 52460 41976
rect 52512 42004 52518 42016
rect 52549 42007 52607 42013
rect 52549 42004 52561 42007
rect 52512 41976 52561 42004
rect 52512 41964 52518 41976
rect 52549 41973 52561 41976
rect 52595 41973 52607 42007
rect 52549 41967 52607 41973
rect 52638 41964 52644 42016
rect 52696 42004 52702 42016
rect 56045 42007 56103 42013
rect 56045 42004 56057 42007
rect 52696 41976 56057 42004
rect 52696 41964 52702 41976
rect 56045 41973 56057 41976
rect 56091 42004 56103 42007
rect 56318 42004 56324 42016
rect 56091 41976 56324 42004
rect 56091 41973 56103 41976
rect 56045 41967 56103 41973
rect 56318 41964 56324 41976
rect 56376 41964 56382 42016
rect 552 41914 66424 41936
rect 552 41862 2918 41914
rect 2970 41862 2982 41914
rect 3034 41862 3046 41914
rect 3098 41862 3110 41914
rect 3162 41862 3174 41914
rect 3226 41862 50918 41914
rect 50970 41862 50982 41914
rect 51034 41862 51046 41914
rect 51098 41862 51110 41914
rect 51162 41862 51174 41914
rect 51226 41862 66424 41914
rect 552 41840 66424 41862
rect 9490 41760 9496 41812
rect 9548 41800 9554 41812
rect 9953 41803 10011 41809
rect 9953 41800 9965 41803
rect 9548 41772 9965 41800
rect 9548 41760 9554 41772
rect 9953 41769 9965 41772
rect 9999 41769 10011 41803
rect 9953 41763 10011 41769
rect 14366 41760 14372 41812
rect 14424 41800 14430 41812
rect 15565 41803 15623 41809
rect 15565 41800 15577 41803
rect 14424 41772 15577 41800
rect 14424 41760 14430 41772
rect 15565 41769 15577 41772
rect 15611 41769 15623 41803
rect 15565 41763 15623 41769
rect 15657 41803 15715 41809
rect 15657 41769 15669 41803
rect 15703 41800 15715 41803
rect 17773 41803 17831 41809
rect 17773 41800 17785 41803
rect 15703 41772 17785 41800
rect 15703 41769 15715 41772
rect 15657 41763 15715 41769
rect 17773 41769 17785 41772
rect 17819 41769 17831 41803
rect 17773 41763 17831 41769
rect 18414 41760 18420 41812
rect 18472 41800 18478 41812
rect 18782 41800 18788 41812
rect 18472 41772 18788 41800
rect 18472 41760 18478 41772
rect 18782 41760 18788 41772
rect 18840 41800 18846 41812
rect 22005 41803 22063 41809
rect 18840 41772 20300 41800
rect 18840 41760 18846 41772
rect 8294 41732 8300 41744
rect 7760 41704 8300 41732
rect 7760 41673 7788 41704
rect 8294 41692 8300 41704
rect 8352 41692 8358 41744
rect 10318 41732 10324 41744
rect 9246 41704 10324 41732
rect 10318 41692 10324 41704
rect 10376 41692 10382 41744
rect 13814 41732 13820 41744
rect 13018 41704 13820 41732
rect 13814 41692 13820 41704
rect 13872 41692 13878 41744
rect 16758 41692 16764 41744
rect 16816 41732 16822 41744
rect 17034 41732 17040 41744
rect 16816 41704 17040 41732
rect 16816 41692 16822 41704
rect 17034 41692 17040 41704
rect 17092 41692 17098 41744
rect 17218 41692 17224 41744
rect 17276 41732 17282 41744
rect 18233 41735 18291 41741
rect 18233 41732 18245 41735
rect 17276 41704 18245 41732
rect 17276 41692 17282 41704
rect 18233 41701 18245 41704
rect 18279 41701 18291 41735
rect 18233 41695 18291 41701
rect 20162 41692 20168 41744
rect 20220 41692 20226 41744
rect 20272 41732 20300 41772
rect 22005 41769 22017 41803
rect 22051 41800 22063 41803
rect 22051 41772 22416 41800
rect 22051 41769 22063 41772
rect 22005 41763 22063 41769
rect 22388 41732 22416 41772
rect 22462 41760 22468 41812
rect 22520 41760 22526 41812
rect 23658 41760 23664 41812
rect 23716 41800 23722 41812
rect 24765 41803 24823 41809
rect 24765 41800 24777 41803
rect 23716 41772 24777 41800
rect 23716 41760 23722 41772
rect 24765 41769 24777 41772
rect 24811 41769 24823 41803
rect 24765 41763 24823 41769
rect 22557 41735 22615 41741
rect 22557 41732 22569 41735
rect 20272 41704 22324 41732
rect 22388 41704 22569 41732
rect 7745 41667 7803 41673
rect 7745 41633 7757 41667
rect 7791 41633 7803 41667
rect 7745 41627 7803 41633
rect 9582 41624 9588 41676
rect 9640 41624 9646 41676
rect 10045 41667 10103 41673
rect 10045 41633 10057 41667
rect 10091 41664 10103 41667
rect 10778 41664 10784 41676
rect 10091 41636 10784 41664
rect 10091 41633 10103 41636
rect 10045 41627 10103 41633
rect 10778 41624 10784 41636
rect 10836 41624 10842 41676
rect 8018 41556 8024 41608
rect 8076 41556 8082 41608
rect 9600 41596 9628 41624
rect 10226 41596 10232 41608
rect 9600 41568 10232 41596
rect 10226 41556 10232 41568
rect 10284 41556 10290 41608
rect 11514 41556 11520 41608
rect 11572 41556 11578 41608
rect 11790 41556 11796 41608
rect 11848 41556 11854 41608
rect 12986 41556 12992 41608
rect 13044 41596 13050 41608
rect 13265 41599 13323 41605
rect 13265 41596 13277 41599
rect 13044 41568 13277 41596
rect 13044 41556 13050 41568
rect 13265 41565 13277 41568
rect 13311 41596 13323 41599
rect 13909 41599 13967 41605
rect 13909 41596 13921 41599
rect 13311 41568 13921 41596
rect 13311 41565 13323 41568
rect 13265 41559 13323 41565
rect 13909 41565 13921 41568
rect 13955 41565 13967 41599
rect 13909 41559 13967 41565
rect 14553 41599 14611 41605
rect 14553 41565 14565 41599
rect 14599 41596 14611 41599
rect 15562 41596 15568 41608
rect 14599 41568 15568 41596
rect 14599 41565 14611 41568
rect 14553 41559 14611 41565
rect 15562 41556 15568 41568
rect 15620 41556 15626 41608
rect 15654 41556 15660 41608
rect 15712 41596 15718 41608
rect 15841 41599 15899 41605
rect 15841 41596 15853 41599
rect 15712 41568 15853 41596
rect 15712 41556 15718 41568
rect 15841 41565 15853 41568
rect 15887 41596 15899 41599
rect 16482 41596 16488 41608
rect 15887 41568 16488 41596
rect 15887 41565 15899 41568
rect 15841 41559 15899 41565
rect 16482 41556 16488 41568
rect 16540 41556 16546 41608
rect 16850 41556 16856 41608
rect 16908 41556 16914 41608
rect 17052 41596 17080 41692
rect 17126 41624 17132 41676
rect 17184 41624 17190 41676
rect 17681 41667 17739 41673
rect 17681 41633 17693 41667
rect 17727 41664 17739 41667
rect 17954 41664 17960 41676
rect 17727 41636 17960 41664
rect 17727 41633 17739 41636
rect 17681 41627 17739 41633
rect 17954 41624 17960 41636
rect 18012 41624 18018 41676
rect 18141 41667 18199 41673
rect 18141 41633 18153 41667
rect 18187 41633 18199 41667
rect 18141 41627 18199 41633
rect 18156 41596 18184 41627
rect 19334 41624 19340 41676
rect 19392 41664 19398 41676
rect 19521 41667 19579 41673
rect 19521 41664 19533 41667
rect 19392 41636 19533 41664
rect 19392 41624 19398 41636
rect 19521 41633 19533 41636
rect 19567 41664 19579 41667
rect 21545 41667 21603 41673
rect 21545 41664 21557 41667
rect 19567 41636 21557 41664
rect 19567 41633 19579 41636
rect 19521 41627 19579 41633
rect 21545 41633 21557 41636
rect 21591 41633 21603 41667
rect 21545 41627 21603 41633
rect 21637 41667 21695 41673
rect 21637 41633 21649 41667
rect 21683 41664 21695 41667
rect 22296 41664 22324 41704
rect 22557 41701 22569 41704
rect 22603 41701 22615 41735
rect 22557 41695 22615 41701
rect 23290 41692 23296 41744
rect 23348 41692 23354 41744
rect 24780 41732 24808 41763
rect 25130 41760 25136 41812
rect 25188 41800 25194 41812
rect 25225 41803 25283 41809
rect 25225 41800 25237 41803
rect 25188 41772 25237 41800
rect 25188 41760 25194 41772
rect 25225 41769 25237 41772
rect 25271 41769 25283 41803
rect 25225 41763 25283 41769
rect 25593 41803 25651 41809
rect 25593 41769 25605 41803
rect 25639 41800 25651 41803
rect 27430 41800 27436 41812
rect 25639 41772 27436 41800
rect 25639 41769 25651 41772
rect 25593 41763 25651 41769
rect 27430 41760 27436 41772
rect 27488 41760 27494 41812
rect 27614 41760 27620 41812
rect 27672 41800 27678 41812
rect 28169 41803 28227 41809
rect 27672 41772 28028 41800
rect 27672 41760 27678 41772
rect 25685 41735 25743 41741
rect 25685 41732 25697 41735
rect 24780 41704 25697 41732
rect 25685 41701 25697 41704
rect 25731 41701 25743 41735
rect 25685 41695 25743 41701
rect 26694 41692 26700 41744
rect 26752 41692 26758 41744
rect 28000 41732 28028 41772
rect 28169 41769 28181 41803
rect 28215 41800 28227 41803
rect 29454 41800 29460 41812
rect 28215 41772 29460 41800
rect 28215 41769 28227 41772
rect 28169 41763 28227 41769
rect 29454 41760 29460 41772
rect 29512 41760 29518 41812
rect 33134 41800 33140 41812
rect 29564 41772 33140 41800
rect 28258 41732 28264 41744
rect 27922 41704 28264 41732
rect 28258 41692 28264 41704
rect 28316 41692 28322 41744
rect 28718 41692 28724 41744
rect 28776 41732 28782 41744
rect 29564 41732 29592 41772
rect 33134 41760 33140 41772
rect 33192 41760 33198 41812
rect 33226 41760 33232 41812
rect 33284 41760 33290 41812
rect 33594 41760 33600 41812
rect 33652 41800 33658 41812
rect 33689 41803 33747 41809
rect 33689 41800 33701 41803
rect 33652 41772 33701 41800
rect 33652 41760 33658 41772
rect 33689 41769 33701 41772
rect 33735 41769 33747 41803
rect 33689 41763 33747 41769
rect 34238 41760 34244 41812
rect 34296 41800 34302 41812
rect 36170 41800 36176 41812
rect 34296 41772 36176 41800
rect 34296 41760 34302 41772
rect 36170 41760 36176 41772
rect 36228 41760 36234 41812
rect 36265 41803 36323 41809
rect 36265 41769 36277 41803
rect 36311 41800 36323 41803
rect 36725 41803 36783 41809
rect 36725 41800 36737 41803
rect 36311 41772 36737 41800
rect 36311 41769 36323 41772
rect 36265 41763 36323 41769
rect 36725 41769 36737 41772
rect 36771 41769 36783 41803
rect 36725 41763 36783 41769
rect 37182 41760 37188 41812
rect 37240 41760 37246 41812
rect 39114 41800 39120 41812
rect 38396 41772 39120 41800
rect 38396 41744 38424 41772
rect 39114 41760 39120 41772
rect 39172 41760 39178 41812
rect 41877 41803 41935 41809
rect 41877 41769 41889 41803
rect 41923 41800 41935 41803
rect 42150 41800 42156 41812
rect 41923 41772 42156 41800
rect 41923 41769 41935 41772
rect 41877 41763 41935 41769
rect 42150 41760 42156 41772
rect 42208 41760 42214 41812
rect 42337 41803 42395 41809
rect 42337 41769 42349 41803
rect 42383 41800 42395 41803
rect 42518 41800 42524 41812
rect 42383 41772 42524 41800
rect 42383 41769 42395 41772
rect 42337 41763 42395 41769
rect 42518 41760 42524 41772
rect 42576 41760 42582 41812
rect 43165 41803 43223 41809
rect 43165 41769 43177 41803
rect 43211 41800 43223 41803
rect 43346 41800 43352 41812
rect 43211 41772 43352 41800
rect 43211 41769 43223 41772
rect 43165 41763 43223 41769
rect 43346 41760 43352 41772
rect 43404 41760 43410 41812
rect 43530 41760 43536 41812
rect 43588 41800 43594 41812
rect 43806 41800 43812 41812
rect 43588 41772 43812 41800
rect 43588 41760 43594 41772
rect 43806 41760 43812 41772
rect 43864 41760 43870 41812
rect 43898 41760 43904 41812
rect 43956 41800 43962 41812
rect 45002 41800 45008 41812
rect 43956 41772 45008 41800
rect 43956 41760 43962 41772
rect 45002 41760 45008 41772
rect 45060 41760 45066 41812
rect 45741 41803 45799 41809
rect 45741 41769 45753 41803
rect 45787 41800 45799 41803
rect 46014 41800 46020 41812
rect 45787 41772 46020 41800
rect 45787 41769 45799 41772
rect 45741 41763 45799 41769
rect 46014 41760 46020 41772
rect 46072 41760 46078 41812
rect 47394 41760 47400 41812
rect 47452 41800 47458 41812
rect 47581 41803 47639 41809
rect 47581 41800 47593 41803
rect 47452 41772 47593 41800
rect 47452 41760 47458 41772
rect 47581 41769 47593 41772
rect 47627 41769 47639 41803
rect 47581 41763 47639 41769
rect 48041 41803 48099 41809
rect 48041 41769 48053 41803
rect 48087 41769 48099 41803
rect 48041 41763 48099 41769
rect 28776 41704 29592 41732
rect 28776 41692 28782 41704
rect 29638 41692 29644 41744
rect 29696 41732 29702 41744
rect 32030 41732 32036 41744
rect 29696 41704 32036 41732
rect 29696 41692 29702 41704
rect 32030 41692 32036 41704
rect 32088 41692 32094 41744
rect 32214 41692 32220 41744
rect 32272 41732 32278 41744
rect 34517 41735 34575 41741
rect 34517 41732 34529 41735
rect 32272 41704 34529 41732
rect 32272 41692 32278 41704
rect 34517 41701 34529 41704
rect 34563 41732 34575 41735
rect 34882 41732 34888 41744
rect 34563 41704 34888 41732
rect 34563 41701 34575 41704
rect 34517 41695 34575 41701
rect 34882 41692 34888 41704
rect 34940 41692 34946 41744
rect 38378 41732 38384 41744
rect 35636 41704 38384 41732
rect 24854 41664 24860 41676
rect 21683 41636 22232 41664
rect 22296 41636 22600 41664
rect 24426 41636 24860 41664
rect 21683 41633 21695 41636
rect 21637 41627 21695 41633
rect 17052 41568 18184 41596
rect 18322 41556 18328 41608
rect 18380 41556 18386 41608
rect 18414 41556 18420 41608
rect 18472 41596 18478 41608
rect 19153 41599 19211 41605
rect 19153 41596 19165 41599
rect 18472 41568 19165 41596
rect 18472 41556 18478 41568
rect 19153 41565 19165 41568
rect 19199 41565 19211 41599
rect 19153 41559 19211 41565
rect 21453 41599 21511 41605
rect 21453 41565 21465 41599
rect 21499 41565 21511 41599
rect 22094 41596 22100 41608
rect 21453 41559 21511 41565
rect 21652 41568 22100 41596
rect 9030 41488 9036 41540
rect 9088 41528 9094 41540
rect 9585 41531 9643 41537
rect 9585 41528 9597 41531
rect 9088 41500 9597 41528
rect 9088 41488 9094 41500
rect 9585 41497 9597 41500
rect 9631 41497 9643 41531
rect 9585 41491 9643 41497
rect 15105 41531 15163 41537
rect 15105 41497 15117 41531
rect 15151 41528 15163 41531
rect 19058 41528 19064 41540
rect 15151 41500 19064 41528
rect 15151 41497 15163 41500
rect 15105 41491 15163 41497
rect 19058 41488 19064 41500
rect 19116 41488 19122 41540
rect 21468 41528 21496 41559
rect 21652 41528 21680 41568
rect 22094 41556 22100 41568
rect 22152 41556 22158 41608
rect 22204 41596 22232 41636
rect 22572 41608 22600 41636
rect 24854 41624 24860 41636
rect 24912 41624 24918 41676
rect 26234 41624 26240 41676
rect 26292 41664 26298 41676
rect 26418 41664 26424 41676
rect 26292 41636 26424 41664
rect 26292 41624 26298 41636
rect 26418 41624 26424 41636
rect 26476 41624 26482 41676
rect 28629 41667 28687 41673
rect 28629 41633 28641 41667
rect 28675 41664 28687 41667
rect 29089 41667 29147 41673
rect 29089 41664 29101 41667
rect 28675 41636 29101 41664
rect 28675 41633 28687 41636
rect 28629 41627 28687 41633
rect 29089 41633 29101 41636
rect 29135 41633 29147 41667
rect 29089 41627 29147 41633
rect 29178 41624 29184 41676
rect 29236 41664 29242 41676
rect 32858 41664 32864 41676
rect 29236 41636 32864 41664
rect 29236 41624 29242 41636
rect 32858 41624 32864 41636
rect 32916 41624 32922 41676
rect 32950 41624 32956 41676
rect 33008 41664 33014 41676
rect 33321 41667 33379 41673
rect 33321 41664 33333 41667
rect 33008 41636 33333 41664
rect 33008 41624 33014 41636
rect 33321 41633 33333 41636
rect 33367 41633 33379 41667
rect 33321 41627 33379 41633
rect 34146 41624 34152 41676
rect 34204 41664 34210 41676
rect 35636 41664 35664 41704
rect 34204 41636 35664 41664
rect 35713 41667 35771 41673
rect 34204 41624 34210 41636
rect 35713 41633 35725 41667
rect 35759 41664 35771 41667
rect 36173 41667 36231 41673
rect 36173 41664 36185 41667
rect 35759 41636 36185 41664
rect 35759 41633 35771 41636
rect 35713 41627 35771 41633
rect 36173 41633 36185 41636
rect 36219 41633 36231 41667
rect 36173 41627 36231 41633
rect 22370 41596 22376 41608
rect 22204 41568 22376 41596
rect 22370 41556 22376 41568
rect 22428 41556 22434 41608
rect 22554 41556 22560 41608
rect 22612 41596 22618 41608
rect 22649 41599 22707 41605
rect 22649 41596 22661 41599
rect 22612 41568 22661 41596
rect 22612 41556 22618 41568
rect 22649 41565 22661 41568
rect 22695 41565 22707 41599
rect 22649 41559 22707 41565
rect 23017 41599 23075 41605
rect 23017 41565 23029 41599
rect 23063 41565 23075 41599
rect 23017 41559 23075 41565
rect 21468 41500 21680 41528
rect 22002 41488 22008 41540
rect 22060 41528 22066 41540
rect 23032 41528 23060 41559
rect 24026 41556 24032 41608
rect 24084 41596 24090 41608
rect 25682 41596 25688 41608
rect 24084 41568 25688 41596
rect 24084 41556 24090 41568
rect 25682 41556 25688 41568
rect 25740 41596 25746 41608
rect 25777 41599 25835 41605
rect 25777 41596 25789 41599
rect 25740 41568 25789 41596
rect 25740 41556 25746 41568
rect 25777 41565 25789 41568
rect 25823 41565 25835 41599
rect 25777 41559 25835 41565
rect 25958 41556 25964 41608
rect 26016 41596 26022 41608
rect 26016 41568 27752 41596
rect 26016 41556 26022 41568
rect 22060 41500 23060 41528
rect 22060 41488 22066 41500
rect 12434 41420 12440 41472
rect 12492 41460 12498 41472
rect 13357 41463 13415 41469
rect 13357 41460 13369 41463
rect 12492 41432 13369 41460
rect 12492 41420 12498 41432
rect 13357 41429 13369 41432
rect 13403 41429 13415 41463
rect 13357 41423 13415 41429
rect 15197 41463 15255 41469
rect 15197 41429 15209 41463
rect 15243 41460 15255 41463
rect 15378 41460 15384 41472
rect 15243 41432 15384 41460
rect 15243 41429 15255 41432
rect 15197 41423 15255 41429
rect 15378 41420 15384 41432
rect 15436 41420 15442 41472
rect 17494 41420 17500 41472
rect 17552 41420 17558 41472
rect 17954 41420 17960 41472
rect 18012 41460 18018 41472
rect 18601 41463 18659 41469
rect 18601 41460 18613 41463
rect 18012 41432 18613 41460
rect 18012 41420 18018 41432
rect 18601 41429 18613 41432
rect 18647 41429 18659 41463
rect 18601 41423 18659 41429
rect 20073 41463 20131 41469
rect 20073 41429 20085 41463
rect 20119 41460 20131 41463
rect 21266 41460 21272 41472
rect 20119 41432 21272 41460
rect 20119 41429 20131 41432
rect 20073 41423 20131 41429
rect 21266 41420 21272 41432
rect 21324 41420 21330 41472
rect 21450 41420 21456 41472
rect 21508 41460 21514 41472
rect 22097 41463 22155 41469
rect 22097 41460 22109 41463
rect 21508 41432 22109 41460
rect 21508 41420 21514 41432
rect 22097 41429 22109 41432
rect 22143 41429 22155 41463
rect 22097 41423 22155 41429
rect 22370 41420 22376 41472
rect 22428 41460 22434 41472
rect 23290 41460 23296 41472
rect 22428 41432 23296 41460
rect 22428 41420 22434 41432
rect 23290 41420 23296 41432
rect 23348 41420 23354 41472
rect 24854 41420 24860 41472
rect 24912 41460 24918 41472
rect 27338 41460 27344 41472
rect 24912 41432 27344 41460
rect 24912 41420 24918 41432
rect 27338 41420 27344 41432
rect 27396 41420 27402 41472
rect 27724 41460 27752 41568
rect 28718 41556 28724 41608
rect 28776 41556 28782 41608
rect 28810 41556 28816 41608
rect 28868 41556 28874 41608
rect 29733 41599 29791 41605
rect 29733 41565 29745 41599
rect 29779 41596 29791 41599
rect 29822 41596 29828 41608
rect 29779 41568 29828 41596
rect 29779 41565 29791 41568
rect 29733 41559 29791 41565
rect 29822 41556 29828 41568
rect 29880 41556 29886 41608
rect 31754 41556 31760 41608
rect 31812 41596 31818 41608
rect 32582 41596 32588 41608
rect 31812 41568 32588 41596
rect 31812 41556 31818 41568
rect 32582 41556 32588 41568
rect 32640 41556 32646 41608
rect 32674 41556 32680 41608
rect 32732 41596 32738 41608
rect 33042 41596 33048 41608
rect 32732 41568 33048 41596
rect 32732 41556 32738 41568
rect 33042 41556 33048 41568
rect 33100 41556 33106 41608
rect 33134 41556 33140 41608
rect 33192 41596 33198 41608
rect 34054 41596 34060 41608
rect 33192 41568 34060 41596
rect 33192 41556 33198 41568
rect 34054 41556 34060 41568
rect 34112 41556 34118 41608
rect 35161 41599 35219 41605
rect 35161 41565 35173 41599
rect 35207 41596 35219 41599
rect 35986 41596 35992 41608
rect 35207 41568 35992 41596
rect 35207 41565 35219 41568
rect 35161 41559 35219 41565
rect 35986 41556 35992 41568
rect 36044 41556 36050 41608
rect 36372 41605 36400 41704
rect 38378 41692 38384 41704
rect 38436 41692 38442 41744
rect 38838 41692 38844 41744
rect 38896 41692 38902 41744
rect 40310 41692 40316 41744
rect 40368 41732 40374 41744
rect 40494 41732 40500 41744
rect 40368 41704 40500 41732
rect 40368 41692 40374 41704
rect 40494 41692 40500 41704
rect 40552 41692 40558 41744
rect 43073 41735 43131 41741
rect 43073 41701 43085 41735
rect 43119 41732 43131 41735
rect 43119 41704 43576 41732
rect 43119 41701 43131 41704
rect 43073 41695 43131 41701
rect 36722 41624 36728 41676
rect 36780 41664 36786 41676
rect 37093 41667 37151 41673
rect 37093 41664 37105 41667
rect 36780 41636 37105 41664
rect 36780 41624 36786 41636
rect 37093 41633 37105 41636
rect 37139 41664 37151 41667
rect 37553 41667 37611 41673
rect 37553 41664 37565 41667
rect 37139 41636 37565 41664
rect 37139 41633 37151 41636
rect 37093 41627 37151 41633
rect 37553 41633 37565 41636
rect 37599 41633 37611 41667
rect 37553 41627 37611 41633
rect 38470 41624 38476 41676
rect 38528 41664 38534 41676
rect 38565 41667 38623 41673
rect 38565 41664 38577 41667
rect 38528 41636 38577 41664
rect 38528 41624 38534 41636
rect 38565 41633 38577 41636
rect 38611 41633 38623 41667
rect 38565 41627 38623 41633
rect 39942 41624 39948 41676
rect 40000 41664 40006 41676
rect 40954 41664 40960 41676
rect 40000 41636 40960 41664
rect 40000 41624 40006 41636
rect 40954 41624 40960 41636
rect 41012 41624 41018 41676
rect 42245 41667 42303 41673
rect 42245 41633 42257 41667
rect 42291 41664 42303 41667
rect 42291 41636 43484 41664
rect 42291 41633 42303 41636
rect 42245 41627 42303 41633
rect 36357 41599 36415 41605
rect 36357 41565 36369 41599
rect 36403 41565 36415 41599
rect 36357 41559 36415 41565
rect 36446 41556 36452 41608
rect 36504 41596 36510 41608
rect 36504 41568 36676 41596
rect 36504 41556 36510 41568
rect 28258 41488 28264 41540
rect 28316 41488 28322 41540
rect 28350 41488 28356 41540
rect 28408 41528 28414 41540
rect 36538 41528 36544 41540
rect 28408 41500 36544 41528
rect 28408 41488 28414 41500
rect 36538 41488 36544 41500
rect 36596 41488 36602 41540
rect 36648 41528 36676 41568
rect 36814 41556 36820 41608
rect 36872 41596 36878 41608
rect 37277 41599 37335 41605
rect 37277 41596 37289 41599
rect 36872 41568 37289 41596
rect 36872 41556 36878 41568
rect 37277 41565 37289 41568
rect 37323 41565 37335 41599
rect 37277 41559 37335 41565
rect 37366 41556 37372 41608
rect 37424 41596 37430 41608
rect 37829 41599 37887 41605
rect 37829 41596 37841 41599
rect 37424 41568 37841 41596
rect 37424 41556 37430 41568
rect 37829 41565 37841 41568
rect 37875 41565 37887 41599
rect 37829 41559 37887 41565
rect 37936 41568 39896 41596
rect 37936 41528 37964 41568
rect 36648 41500 37964 41528
rect 30374 41460 30380 41472
rect 27724 41432 30380 41460
rect 30374 41420 30380 41432
rect 30432 41420 30438 41472
rect 35802 41420 35808 41472
rect 35860 41420 35866 41472
rect 35986 41420 35992 41472
rect 36044 41460 36050 41472
rect 36630 41460 36636 41472
rect 36044 41432 36636 41460
rect 36044 41420 36050 41432
rect 36630 41420 36636 41432
rect 36688 41420 36694 41472
rect 38473 41463 38531 41469
rect 38473 41429 38485 41463
rect 38519 41460 38531 41463
rect 38930 41460 38936 41472
rect 38519 41432 38936 41460
rect 38519 41429 38531 41432
rect 38473 41423 38531 41429
rect 38930 41420 38936 41432
rect 38988 41420 38994 41472
rect 39868 41460 39896 41568
rect 40218 41556 40224 41608
rect 40276 41596 40282 41608
rect 40313 41599 40371 41605
rect 40313 41596 40325 41599
rect 40276 41568 40325 41596
rect 40276 41556 40282 41568
rect 40313 41565 40325 41568
rect 40359 41565 40371 41599
rect 40313 41559 40371 41565
rect 41782 41556 41788 41608
rect 41840 41596 41846 41608
rect 42518 41596 42524 41608
rect 41840 41568 42524 41596
rect 41840 41556 41846 41568
rect 42518 41556 42524 41568
rect 42576 41556 42582 41608
rect 43162 41596 43168 41608
rect 43088 41568 43168 41596
rect 40770 41488 40776 41540
rect 40828 41528 40834 41540
rect 43088 41528 43116 41568
rect 43162 41556 43168 41568
rect 43220 41596 43226 41608
rect 43349 41599 43407 41605
rect 43349 41596 43361 41599
rect 43220 41568 43361 41596
rect 43220 41556 43226 41568
rect 43349 41565 43361 41568
rect 43395 41565 43407 41599
rect 43349 41559 43407 41565
rect 40828 41500 43116 41528
rect 43456 41528 43484 41636
rect 43548 41596 43576 41704
rect 43622 41692 43628 41744
rect 43680 41732 43686 41744
rect 44177 41735 44235 41741
rect 44177 41732 44189 41735
rect 43680 41704 44189 41732
rect 43680 41692 43686 41704
rect 44177 41701 44189 41704
rect 44223 41732 44235 41735
rect 44223 41704 45140 41732
rect 44223 41701 44235 41704
rect 44177 41695 44235 41701
rect 43806 41624 43812 41676
rect 43864 41664 43870 41676
rect 44085 41667 44143 41673
rect 44085 41664 44097 41667
rect 43864 41636 44097 41664
rect 43864 41624 43870 41636
rect 44085 41633 44097 41636
rect 44131 41633 44143 41667
rect 44726 41664 44732 41676
rect 44085 41627 44143 41633
rect 44284 41636 44732 41664
rect 44284 41596 44312 41636
rect 44726 41624 44732 41636
rect 44784 41624 44790 41676
rect 45112 41673 45140 41704
rect 45922 41692 45928 41744
rect 45980 41732 45986 41744
rect 46109 41735 46167 41741
rect 46109 41732 46121 41735
rect 45980 41704 46121 41732
rect 45980 41692 45986 41704
rect 46109 41701 46121 41704
rect 46155 41701 46167 41735
rect 46109 41695 46167 41701
rect 46750 41692 46756 41744
rect 46808 41732 46814 41744
rect 48056 41732 48084 41763
rect 48130 41760 48136 41812
rect 48188 41760 48194 41812
rect 48498 41760 48504 41812
rect 48556 41760 48562 41812
rect 50430 41800 50436 41812
rect 49712 41772 50436 41800
rect 49712 41741 49740 41772
rect 50430 41760 50436 41772
rect 50488 41760 50494 41812
rect 52362 41760 52368 41812
rect 52420 41800 52426 41812
rect 53009 41803 53067 41809
rect 53009 41800 53021 41803
rect 52420 41772 53021 41800
rect 52420 41760 52426 41772
rect 53009 41769 53021 41772
rect 53055 41769 53067 41803
rect 53009 41763 53067 41769
rect 48593 41735 48651 41741
rect 48593 41732 48605 41735
rect 46808 41704 47979 41732
rect 48056 41704 48605 41732
rect 46808 41692 46814 41704
rect 45097 41667 45155 41673
rect 45097 41633 45109 41667
rect 45143 41633 45155 41667
rect 45097 41627 45155 41633
rect 47673 41667 47731 41673
rect 47673 41633 47685 41667
rect 47719 41664 47731 41667
rect 47854 41664 47860 41676
rect 47719 41636 47860 41664
rect 47719 41633 47731 41636
rect 47673 41627 47731 41633
rect 47854 41624 47860 41636
rect 47912 41624 47918 41676
rect 43548 41568 44312 41596
rect 44361 41599 44419 41605
rect 44361 41565 44373 41599
rect 44407 41596 44419 41599
rect 44407 41568 44680 41596
rect 44407 41565 44419 41568
rect 44361 41559 44419 41565
rect 44545 41531 44603 41537
rect 44545 41528 44557 41531
rect 43456 41500 44557 41528
rect 40828 41488 40834 41500
rect 44545 41497 44557 41500
rect 44591 41497 44603 41531
rect 44545 41491 44603 41497
rect 40678 41460 40684 41472
rect 39868 41432 40684 41460
rect 40678 41420 40684 41432
rect 40736 41420 40742 41472
rect 42702 41420 42708 41472
rect 42760 41420 42766 41472
rect 43254 41420 43260 41472
rect 43312 41460 43318 41472
rect 43717 41463 43775 41469
rect 43717 41460 43729 41463
rect 43312 41432 43729 41460
rect 43312 41420 43318 41432
rect 43717 41429 43729 41432
rect 43763 41429 43775 41463
rect 43717 41423 43775 41429
rect 43806 41420 43812 41472
rect 43864 41460 43870 41472
rect 44082 41460 44088 41472
rect 43864 41432 44088 41460
rect 43864 41420 43870 41432
rect 44082 41420 44088 41432
rect 44140 41460 44146 41472
rect 44652 41460 44680 41568
rect 45830 41556 45836 41608
rect 45888 41596 45894 41608
rect 46201 41599 46259 41605
rect 46201 41596 46213 41599
rect 45888 41568 46213 41596
rect 45888 41556 45894 41568
rect 46201 41565 46213 41568
rect 46247 41565 46259 41599
rect 46201 41559 46259 41565
rect 46385 41599 46443 41605
rect 46385 41565 46397 41599
rect 46431 41596 46443 41599
rect 46842 41596 46848 41608
rect 46431 41568 46848 41596
rect 46431 41565 46443 41568
rect 46385 41559 46443 41565
rect 45738 41488 45744 41540
rect 45796 41528 45802 41540
rect 45922 41528 45928 41540
rect 45796 41500 45928 41528
rect 45796 41488 45802 41500
rect 45922 41488 45928 41500
rect 45980 41528 45986 41540
rect 46400 41528 46428 41559
rect 46842 41556 46848 41568
rect 46900 41596 46906 41608
rect 47397 41599 47455 41605
rect 47397 41596 47409 41599
rect 46900 41568 47409 41596
rect 46900 41556 46906 41568
rect 47397 41565 47409 41568
rect 47443 41596 47455 41599
rect 47578 41596 47584 41608
rect 47443 41568 47584 41596
rect 47443 41565 47455 41568
rect 47397 41559 47455 41565
rect 47578 41556 47584 41568
rect 47636 41556 47642 41608
rect 47951 41596 47979 41704
rect 48593 41701 48605 41704
rect 48639 41701 48651 41735
rect 48593 41695 48651 41701
rect 49697 41735 49755 41741
rect 49697 41701 49709 41735
rect 49743 41701 49755 41735
rect 49697 41695 49755 41701
rect 50338 41692 50344 41744
rect 50396 41692 50402 41744
rect 52549 41667 52607 41673
rect 52549 41633 52561 41667
rect 52595 41664 52607 41667
rect 53745 41667 53803 41673
rect 53745 41664 53757 41667
rect 52595 41636 53757 41664
rect 52595 41633 52607 41636
rect 52549 41627 52607 41633
rect 53745 41633 53757 41636
rect 53791 41633 53803 41667
rect 53745 41627 53803 41633
rect 55217 41667 55275 41673
rect 55217 41633 55229 41667
rect 55263 41664 55275 41667
rect 55953 41667 56011 41673
rect 55953 41664 55965 41667
rect 55263 41636 55965 41664
rect 55263 41633 55275 41636
rect 55217 41627 55275 41633
rect 55953 41633 55965 41636
rect 55999 41633 56011 41667
rect 55953 41627 56011 41633
rect 48406 41596 48412 41608
rect 47951 41568 48412 41596
rect 48406 41556 48412 41568
rect 48464 41596 48470 41608
rect 48685 41599 48743 41605
rect 48685 41596 48697 41599
rect 48464 41568 48697 41596
rect 48464 41556 48470 41568
rect 48685 41565 48697 41568
rect 48731 41596 48743 41599
rect 49142 41596 49148 41608
rect 48731 41568 49148 41596
rect 48731 41565 48743 41568
rect 48685 41559 48743 41565
rect 49142 41556 49148 41568
rect 49200 41556 49206 41608
rect 49421 41599 49479 41605
rect 49421 41565 49433 41599
rect 49467 41565 49479 41599
rect 49421 41559 49479 41565
rect 45980 41500 46428 41528
rect 45980 41488 45986 41500
rect 46934 41488 46940 41540
rect 46992 41528 46998 41540
rect 48130 41528 48136 41540
rect 46992 41500 48136 41528
rect 46992 41488 46998 41500
rect 48130 41488 48136 41500
rect 48188 41528 48194 41540
rect 49436 41528 49464 41559
rect 50706 41556 50712 41608
rect 50764 41596 50770 41608
rect 51445 41599 51503 41605
rect 51445 41596 51457 41599
rect 50764 41568 51457 41596
rect 50764 41556 50770 41568
rect 51445 41565 51457 41568
rect 51491 41565 51503 41599
rect 51445 41559 51503 41565
rect 52362 41556 52368 41608
rect 52420 41596 52426 41608
rect 52641 41599 52699 41605
rect 52641 41596 52653 41599
rect 52420 41568 52653 41596
rect 52420 41556 52426 41568
rect 52641 41565 52653 41568
rect 52687 41565 52699 41599
rect 52641 41559 52699 41565
rect 52825 41599 52883 41605
rect 52825 41565 52837 41599
rect 52871 41596 52883 41599
rect 52914 41596 52920 41608
rect 52871 41568 52920 41596
rect 52871 41565 52883 41568
rect 52825 41559 52883 41565
rect 52914 41556 52920 41568
rect 52972 41556 52978 41608
rect 53653 41599 53711 41605
rect 53653 41565 53665 41599
rect 53699 41565 53711 41599
rect 53653 41559 53711 41565
rect 48188 41500 49464 41528
rect 48188 41488 48194 41500
rect 51350 41488 51356 41540
rect 51408 41528 51414 41540
rect 53668 41528 53696 41559
rect 53834 41556 53840 41608
rect 53892 41596 53898 41608
rect 54297 41599 54355 41605
rect 54297 41596 54309 41599
rect 53892 41568 54309 41596
rect 53892 41556 53898 41568
rect 54297 41565 54309 41568
rect 54343 41565 54355 41599
rect 54297 41559 54355 41565
rect 55306 41556 55312 41608
rect 55364 41556 55370 41608
rect 55493 41599 55551 41605
rect 55493 41565 55505 41599
rect 55539 41565 55551 41599
rect 55493 41559 55551 41565
rect 55508 41528 55536 41559
rect 56502 41556 56508 41608
rect 56560 41596 56566 41608
rect 56597 41599 56655 41605
rect 56597 41596 56609 41599
rect 56560 41568 56609 41596
rect 56560 41556 56566 41568
rect 56597 41565 56609 41568
rect 56643 41565 56655 41599
rect 56597 41559 56655 41565
rect 57422 41528 57428 41540
rect 51408 41500 53696 41528
rect 53760 41500 57428 41528
rect 51408 41488 51414 41500
rect 44140 41432 44680 41460
rect 52181 41463 52239 41469
rect 44140 41420 44146 41432
rect 52181 41429 52193 41463
rect 52227 41460 52239 41463
rect 52454 41460 52460 41472
rect 52227 41432 52460 41460
rect 52227 41429 52239 41432
rect 52181 41423 52239 41429
rect 52454 41420 52460 41432
rect 52512 41420 52518 41472
rect 52546 41420 52552 41472
rect 52604 41460 52610 41472
rect 52822 41460 52828 41472
rect 52604 41432 52828 41460
rect 52604 41420 52610 41432
rect 52822 41420 52828 41432
rect 52880 41420 52886 41472
rect 52914 41420 52920 41472
rect 52972 41460 52978 41472
rect 53760 41460 53788 41500
rect 57422 41488 57428 41500
rect 57480 41488 57486 41540
rect 52972 41432 53788 41460
rect 54849 41463 54907 41469
rect 52972 41420 52978 41432
rect 54849 41429 54861 41463
rect 54895 41460 54907 41463
rect 55030 41460 55036 41472
rect 54895 41432 55036 41460
rect 54895 41429 54907 41432
rect 54849 41423 54907 41429
rect 55030 41420 55036 41432
rect 55088 41420 55094 41472
rect 552 41370 66424 41392
rect 552 41318 1998 41370
rect 2050 41318 2062 41370
rect 2114 41318 2126 41370
rect 2178 41318 2190 41370
rect 2242 41318 2254 41370
rect 2306 41318 49998 41370
rect 50050 41318 50062 41370
rect 50114 41318 50126 41370
rect 50178 41318 50190 41370
rect 50242 41318 50254 41370
rect 50306 41318 66424 41370
rect 552 41296 66424 41318
rect 9674 41216 9680 41268
rect 9732 41256 9738 41268
rect 10137 41259 10195 41265
rect 10137 41256 10149 41259
rect 9732 41228 10149 41256
rect 9732 41216 9738 41228
rect 10137 41225 10149 41228
rect 10183 41225 10195 41259
rect 10137 41219 10195 41225
rect 7653 41123 7711 41129
rect 7653 41089 7665 41123
rect 7699 41120 7711 41123
rect 8294 41120 8300 41132
rect 7699 41092 8300 41120
rect 7699 41089 7711 41092
rect 7653 41083 7711 41089
rect 8294 41080 8300 41092
rect 8352 41080 8358 41132
rect 8386 41080 8392 41132
rect 8444 41080 8450 41132
rect 10152 41052 10180 41219
rect 11790 41216 11796 41268
rect 11848 41216 11854 41268
rect 12066 41216 12072 41268
rect 12124 41256 12130 41268
rect 13262 41256 13268 41268
rect 12124 41228 13268 41256
rect 12124 41216 12130 41228
rect 13262 41216 13268 41228
rect 13320 41216 13326 41268
rect 15838 41216 15844 41268
rect 15896 41256 15902 41268
rect 16482 41256 16488 41268
rect 15896 41228 16488 41256
rect 15896 41216 15902 41228
rect 16482 41216 16488 41228
rect 16540 41216 16546 41268
rect 16758 41216 16764 41268
rect 16816 41216 16822 41268
rect 17126 41216 17132 41268
rect 17184 41256 17190 41268
rect 17862 41256 17868 41268
rect 17184 41228 17868 41256
rect 17184 41216 17190 41228
rect 17862 41216 17868 41228
rect 17920 41216 17926 41268
rect 20272 41228 26924 41256
rect 10226 41148 10232 41200
rect 10284 41188 10290 41200
rect 12618 41188 12624 41200
rect 10284 41160 12624 41188
rect 10284 41148 10290 41160
rect 10888 41129 10916 41160
rect 12618 41148 12624 41160
rect 12676 41188 12682 41200
rect 12676 41160 12940 41188
rect 12676 41148 12682 41160
rect 12912 41132 12940 41160
rect 13722 41148 13728 41200
rect 13780 41188 13786 41200
rect 13780 41160 14228 41188
rect 13780 41148 13786 41160
rect 10873 41123 10931 41129
rect 10873 41089 10885 41123
rect 10919 41089 10931 41123
rect 10873 41083 10931 41089
rect 11606 41080 11612 41132
rect 11664 41120 11670 41132
rect 12345 41123 12403 41129
rect 12345 41120 12357 41123
rect 11664 41092 12357 41120
rect 11664 41080 11670 41092
rect 12345 41089 12357 41092
rect 12391 41089 12403 41123
rect 12345 41083 12403 41089
rect 12894 41080 12900 41132
rect 12952 41120 12958 41132
rect 13173 41123 13231 41129
rect 13173 41120 13185 41123
rect 12952 41092 13185 41120
rect 12952 41080 12958 41092
rect 13173 41089 13185 41092
rect 13219 41089 13231 41123
rect 13173 41083 13231 41089
rect 13262 41080 13268 41132
rect 13320 41120 13326 41132
rect 14093 41123 14151 41129
rect 14093 41120 14105 41123
rect 13320 41092 14105 41120
rect 13320 41080 13326 41092
rect 14093 41089 14105 41092
rect 14139 41089 14151 41123
rect 14200 41120 14228 41160
rect 16850 41148 16856 41200
rect 16908 41188 16914 41200
rect 17586 41188 17592 41200
rect 16908 41160 17592 41188
rect 16908 41148 16914 41160
rect 17586 41148 17592 41160
rect 17644 41188 17650 41200
rect 17644 41160 18092 41188
rect 17644 41148 17650 41160
rect 18064 41129 18092 41160
rect 18708 41160 19380 41188
rect 17865 41123 17923 41129
rect 17865 41120 17877 41123
rect 14200 41092 17877 41120
rect 14093 41083 14151 41089
rect 17865 41089 17877 41092
rect 17911 41089 17923 41123
rect 17865 41083 17923 41089
rect 18049 41123 18107 41129
rect 18049 41089 18061 41123
rect 18095 41120 18107 41123
rect 18598 41120 18604 41132
rect 18095 41092 18604 41120
rect 18095 41089 18107 41092
rect 18049 41083 18107 41089
rect 18598 41080 18604 41092
rect 18656 41080 18662 41132
rect 10597 41055 10655 41061
rect 10597 41052 10609 41055
rect 10152 41024 10609 41052
rect 10597 41021 10609 41024
rect 10643 41021 10655 41055
rect 10597 41015 10655 41021
rect 12161 41055 12219 41061
rect 12161 41021 12173 41055
rect 12207 41052 12219 41055
rect 12434 41052 12440 41064
rect 12207 41024 12440 41052
rect 12207 41021 12219 41024
rect 12161 41015 12219 41021
rect 12434 41012 12440 41024
rect 12492 41012 12498 41064
rect 12986 41012 12992 41064
rect 13044 41012 13050 41064
rect 13081 41055 13139 41061
rect 13081 41021 13093 41055
rect 13127 41052 13139 41055
rect 13127 41024 13676 41052
rect 13127 41021 13139 41024
rect 13081 41015 13139 41021
rect 7837 40987 7895 40993
rect 7837 40953 7849 40987
rect 7883 40984 7895 40987
rect 8570 40984 8576 40996
rect 7883 40956 8576 40984
rect 7883 40953 7895 40956
rect 7837 40947 7895 40953
rect 8570 40944 8576 40956
rect 8628 40944 8634 40996
rect 8665 40987 8723 40993
rect 8665 40953 8677 40987
rect 8711 40953 8723 40987
rect 10318 40984 10324 40996
rect 9890 40956 10324 40984
rect 8665 40947 8723 40953
rect 7742 40876 7748 40928
rect 7800 40876 7806 40928
rect 8205 40919 8263 40925
rect 8205 40885 8217 40919
rect 8251 40916 8263 40919
rect 8680 40916 8708 40947
rect 10318 40944 10324 40956
rect 10376 40944 10382 40996
rect 12253 40987 12311 40993
rect 12253 40953 12265 40987
rect 12299 40984 12311 40987
rect 12299 40956 13584 40984
rect 12299 40953 12311 40956
rect 12253 40947 12311 40953
rect 8251 40888 8708 40916
rect 8251 40885 8263 40888
rect 8205 40879 8263 40885
rect 10226 40876 10232 40928
rect 10284 40876 10290 40928
rect 10689 40919 10747 40925
rect 10689 40885 10701 40919
rect 10735 40916 10747 40919
rect 11330 40916 11336 40928
rect 10735 40888 11336 40916
rect 10735 40885 10747 40888
rect 10689 40879 10747 40885
rect 11330 40876 11336 40888
rect 11388 40876 11394 40928
rect 12434 40876 12440 40928
rect 12492 40916 12498 40928
rect 13556 40925 13584 40956
rect 12621 40919 12679 40925
rect 12621 40916 12633 40919
rect 12492 40888 12633 40916
rect 12492 40876 12498 40888
rect 12621 40885 12633 40888
rect 12667 40885 12679 40919
rect 12621 40879 12679 40885
rect 13541 40919 13599 40925
rect 13541 40885 13553 40919
rect 13587 40885 13599 40919
rect 13648 40916 13676 41024
rect 13814 41012 13820 41064
rect 13872 41052 13878 41064
rect 15010 41052 15016 41064
rect 13872 41024 15016 41052
rect 13872 41012 13878 41024
rect 15010 41012 15016 41024
rect 15068 41012 15074 41064
rect 17313 41055 17371 41061
rect 17313 41021 17325 41055
rect 17359 41052 17371 41055
rect 17773 41055 17831 41061
rect 17773 41052 17785 41055
rect 17359 41024 17785 41052
rect 17359 41021 17371 41024
rect 17313 41015 17371 41021
rect 17773 41021 17785 41024
rect 17819 41052 17831 41055
rect 18708 41052 18736 41160
rect 18782 41080 18788 41132
rect 18840 41120 18846 41132
rect 19245 41123 19303 41129
rect 19245 41120 19257 41123
rect 18840 41092 19257 41120
rect 18840 41080 18846 41092
rect 19245 41089 19257 41092
rect 19291 41089 19303 41123
rect 19352 41120 19380 41160
rect 20162 41148 20168 41200
rect 20220 41148 20226 41200
rect 20272 41120 20300 41228
rect 19352 41092 20300 41120
rect 21560 41160 21772 41188
rect 19245 41083 19303 41089
rect 17819 41024 18736 41052
rect 17819 41021 17831 41024
rect 17773 41015 17831 41021
rect 19058 41012 19064 41064
rect 19116 41012 19122 41064
rect 13998 40944 14004 40996
rect 14056 40944 14062 40996
rect 15194 40944 15200 40996
rect 15252 40984 15258 40996
rect 15289 40987 15347 40993
rect 15289 40984 15301 40987
rect 15252 40956 15301 40984
rect 15252 40944 15258 40956
rect 15289 40953 15301 40956
rect 15335 40953 15347 40987
rect 15289 40947 15347 40953
rect 15746 40944 15752 40996
rect 15804 40944 15810 40996
rect 17494 40944 17500 40996
rect 17552 40984 17558 40996
rect 19153 40987 19211 40993
rect 19153 40984 19165 40987
rect 17552 40956 19165 40984
rect 17552 40944 17558 40956
rect 19153 40953 19165 40956
rect 19199 40953 19211 40987
rect 19153 40947 19211 40953
rect 19518 40944 19524 40996
rect 19576 40984 19582 40996
rect 21560 40984 21588 41160
rect 21744 41120 21772 41160
rect 23290 41148 23296 41200
rect 23348 41188 23354 41200
rect 23477 41191 23535 41197
rect 23477 41188 23489 41191
rect 23348 41160 23489 41188
rect 23348 41148 23354 41160
rect 23477 41157 23489 41160
rect 23523 41188 23535 41191
rect 23750 41188 23756 41200
rect 23523 41160 23756 41188
rect 23523 41157 23535 41160
rect 23477 41151 23535 41157
rect 23750 41148 23756 41160
rect 23808 41148 23814 41200
rect 26786 41188 26792 41200
rect 24228 41160 26792 41188
rect 21744 41092 24164 41120
rect 21729 41055 21787 41061
rect 21729 41021 21741 41055
rect 21775 41021 21787 41055
rect 21729 41015 21787 41021
rect 21637 40987 21695 40993
rect 21637 40984 21649 40987
rect 19576 40956 21649 40984
rect 19576 40944 19582 40956
rect 21637 40953 21649 40956
rect 21683 40953 21695 40987
rect 21637 40947 21695 40953
rect 13906 40916 13912 40928
rect 13648 40888 13912 40916
rect 13541 40879 13599 40885
rect 13906 40876 13912 40888
rect 13964 40876 13970 40928
rect 14550 40876 14556 40928
rect 14608 40916 14614 40928
rect 17126 40916 17132 40928
rect 14608 40888 17132 40916
rect 14608 40876 14614 40888
rect 17126 40876 17132 40888
rect 17184 40876 17190 40928
rect 17402 40876 17408 40928
rect 17460 40876 17466 40928
rect 18690 40876 18696 40928
rect 18748 40876 18754 40928
rect 20162 40876 20168 40928
rect 20220 40916 20226 40928
rect 21744 40916 21772 41015
rect 22002 40944 22008 40996
rect 22060 40944 22066 40996
rect 23014 40944 23020 40996
rect 23072 40944 23078 40996
rect 24136 40984 24164 41092
rect 24228 41061 24256 41160
rect 26786 41148 26792 41160
rect 26844 41148 26850 41200
rect 26896 41188 26924 41228
rect 27982 41216 27988 41268
rect 28040 41256 28046 41268
rect 28997 41259 29055 41265
rect 28997 41256 29009 41259
rect 28040 41228 29009 41256
rect 28040 41216 28046 41228
rect 28997 41225 29009 41228
rect 29043 41225 29055 41259
rect 28997 41219 29055 41225
rect 30374 41216 30380 41268
rect 30432 41256 30438 41268
rect 30432 41228 32904 41256
rect 30432 41216 30438 41228
rect 32876 41188 32904 41228
rect 32950 41216 32956 41268
rect 33008 41216 33014 41268
rect 34790 41216 34796 41268
rect 34848 41256 34854 41268
rect 36906 41256 36912 41268
rect 34848 41228 36912 41256
rect 34848 41216 34854 41228
rect 36906 41216 36912 41228
rect 36964 41256 36970 41268
rect 43438 41256 43444 41268
rect 36964 41228 43444 41256
rect 36964 41216 36970 41228
rect 43438 41216 43444 41228
rect 43496 41256 43502 41268
rect 43496 41228 51074 41256
rect 43496 41216 43502 41228
rect 34698 41188 34704 41200
rect 26896 41160 31754 41188
rect 32876 41160 34704 41188
rect 24486 41080 24492 41132
rect 24544 41080 24550 41132
rect 26602 41080 26608 41132
rect 26660 41080 26666 41132
rect 28902 41080 28908 41132
rect 28960 41120 28966 41132
rect 29641 41123 29699 41129
rect 29641 41120 29653 41123
rect 28960 41092 29653 41120
rect 28960 41080 28966 41092
rect 29641 41089 29653 41092
rect 29687 41120 29699 41123
rect 30006 41120 30012 41132
rect 29687 41092 30012 41120
rect 29687 41089 29699 41092
rect 29641 41083 29699 41089
rect 30006 41080 30012 41092
rect 30064 41080 30070 41132
rect 30926 41120 30932 41132
rect 30300 41092 30932 41120
rect 24213 41055 24271 41061
rect 24213 41021 24225 41055
rect 24259 41021 24271 41055
rect 28261 41055 28319 41061
rect 28261 41052 28273 41055
rect 24213 41015 24271 41021
rect 24596 41024 28273 41052
rect 24596 40984 24624 41024
rect 28261 41021 28273 41024
rect 28307 41052 28319 41055
rect 28350 41052 28356 41064
rect 28307 41024 28356 41052
rect 28307 41021 28319 41024
rect 28261 41015 28319 41021
rect 28350 41012 28356 41024
rect 28408 41012 28414 41064
rect 29365 41055 29423 41061
rect 29365 41021 29377 41055
rect 29411 41052 29423 41055
rect 30300 41052 30328 41092
rect 30926 41080 30932 41092
rect 30984 41080 30990 41132
rect 31726 41120 31754 41160
rect 34698 41148 34704 41160
rect 34756 41148 34762 41200
rect 36630 41148 36636 41200
rect 36688 41148 36694 41200
rect 40034 41188 40040 41200
rect 39776 41160 40040 41188
rect 33226 41120 33232 41132
rect 31726 41092 33232 41120
rect 33226 41080 33232 41092
rect 33284 41080 33290 41132
rect 33410 41080 33416 41132
rect 33468 41120 33474 41132
rect 33781 41123 33839 41129
rect 33781 41120 33793 41123
rect 33468 41092 33793 41120
rect 33468 41080 33474 41092
rect 33781 41089 33793 41092
rect 33827 41120 33839 41123
rect 34146 41120 34152 41132
rect 33827 41092 34152 41120
rect 33827 41089 33839 41092
rect 33781 41083 33839 41089
rect 34146 41080 34152 41092
rect 34204 41080 34210 41132
rect 34885 41123 34943 41129
rect 34885 41089 34897 41123
rect 34931 41120 34943 41123
rect 35618 41120 35624 41132
rect 34931 41092 35624 41120
rect 34931 41089 34943 41092
rect 34885 41083 34943 41089
rect 35618 41080 35624 41092
rect 35676 41080 35682 41132
rect 36722 41080 36728 41132
rect 36780 41080 36786 41132
rect 37921 41123 37979 41129
rect 37921 41089 37933 41123
rect 37967 41120 37979 41123
rect 38102 41120 38108 41132
rect 37967 41092 38108 41120
rect 37967 41089 37979 41092
rect 37921 41083 37979 41089
rect 38102 41080 38108 41092
rect 38160 41120 38166 41132
rect 38657 41123 38715 41129
rect 38657 41120 38669 41123
rect 38160 41092 38669 41120
rect 38160 41080 38166 41092
rect 38657 41089 38669 41092
rect 38703 41089 38715 41123
rect 38657 41083 38715 41089
rect 39574 41080 39580 41132
rect 39632 41120 39638 41132
rect 39776 41129 39804 41160
rect 40034 41148 40040 41160
rect 40092 41148 40098 41200
rect 44082 41148 44088 41200
rect 44140 41188 44146 41200
rect 44453 41191 44511 41197
rect 44453 41188 44465 41191
rect 44140 41160 44465 41188
rect 44140 41148 44146 41160
rect 44453 41157 44465 41160
rect 44499 41157 44511 41191
rect 44453 41151 44511 41157
rect 44726 41148 44732 41200
rect 44784 41188 44790 41200
rect 46201 41191 46259 41197
rect 46201 41188 46213 41191
rect 44784 41160 46213 41188
rect 44784 41148 44790 41160
rect 46201 41157 46213 41160
rect 46247 41157 46259 41191
rect 46201 41151 46259 41157
rect 48498 41148 48504 41200
rect 48556 41188 48562 41200
rect 49510 41188 49516 41200
rect 48556 41160 49516 41188
rect 48556 41148 48562 41160
rect 49510 41148 49516 41160
rect 49568 41148 49574 41200
rect 39761 41123 39819 41129
rect 39761 41120 39773 41123
rect 39632 41092 39773 41120
rect 39632 41080 39638 41092
rect 39761 41089 39773 41092
rect 39807 41089 39819 41123
rect 39761 41083 39819 41089
rect 39945 41123 40003 41129
rect 39945 41089 39957 41123
rect 39991 41120 40003 41123
rect 40126 41120 40132 41132
rect 39991 41092 40132 41120
rect 39991 41089 40003 41092
rect 39945 41083 40003 41089
rect 40126 41080 40132 41092
rect 40184 41080 40190 41132
rect 40494 41080 40500 41132
rect 40552 41120 40558 41132
rect 41690 41120 41696 41132
rect 40552 41092 41696 41120
rect 40552 41080 40558 41092
rect 41690 41080 41696 41092
rect 41748 41120 41754 41132
rect 42429 41123 42487 41129
rect 42429 41120 42441 41123
rect 41748 41092 42441 41120
rect 41748 41080 41754 41092
rect 42429 41089 42441 41092
rect 42475 41089 42487 41123
rect 42429 41083 42487 41089
rect 44177 41123 44235 41129
rect 44177 41089 44189 41123
rect 44223 41089 44235 41123
rect 44177 41083 44235 41089
rect 29411 41024 30328 41052
rect 30469 41055 30527 41061
rect 29411 41021 29423 41024
rect 29365 41015 29423 41021
rect 30469 41021 30481 41055
rect 30515 41052 30527 41055
rect 30558 41052 30564 41064
rect 30515 41024 30564 41052
rect 30515 41021 30527 41024
rect 30469 41015 30527 41021
rect 30558 41012 30564 41024
rect 30616 41012 30622 41064
rect 31478 41012 31484 41064
rect 31536 41052 31542 41064
rect 31849 41055 31907 41061
rect 31849 41052 31861 41055
rect 31536 41024 31861 41052
rect 31536 41012 31542 41024
rect 31849 41021 31861 41024
rect 31895 41021 31907 41055
rect 31849 41015 31907 41021
rect 32309 41055 32367 41061
rect 32309 41021 32321 41055
rect 32355 41052 32367 41055
rect 32355 41024 33640 41052
rect 32355 41021 32367 41024
rect 32309 41015 32367 41021
rect 24136 40956 24624 40984
rect 24670 40944 24676 40996
rect 24728 40944 24734 40996
rect 24762 40944 24768 40996
rect 24820 40984 24826 40996
rect 32766 40984 32772 40996
rect 24820 40956 32772 40984
rect 24820 40944 24826 40956
rect 32766 40944 32772 40956
rect 32824 40944 32830 40996
rect 32861 40987 32919 40993
rect 32861 40953 32873 40987
rect 32907 40984 32919 40987
rect 33505 40987 33563 40993
rect 33505 40984 33517 40987
rect 32907 40956 33517 40984
rect 32907 40953 32919 40956
rect 32861 40947 32919 40953
rect 33505 40953 33517 40956
rect 33551 40953 33563 40987
rect 33612 40984 33640 41024
rect 33686 41012 33692 41064
rect 33744 41052 33750 41064
rect 34701 41055 34759 41061
rect 34701 41052 34713 41055
rect 33744 41024 34713 41052
rect 33744 41012 33750 41024
rect 34701 41021 34713 41024
rect 34747 41021 34759 41055
rect 34701 41015 34759 41021
rect 36170 41012 36176 41064
rect 36228 41052 36234 41064
rect 36228 41024 36294 41052
rect 36228 41012 36234 41024
rect 37642 41012 37648 41064
rect 37700 41052 37706 41064
rect 37737 41055 37795 41061
rect 37737 41052 37749 41055
rect 37700 41024 37749 41052
rect 37700 41012 37706 41024
rect 37737 41021 37749 41024
rect 37783 41021 37795 41055
rect 37737 41015 37795 41021
rect 38470 41012 38476 41064
rect 38528 41052 38534 41064
rect 42242 41052 42248 41064
rect 38528 41024 42248 41052
rect 38528 41012 38534 41024
rect 42242 41012 42248 41024
rect 42300 41012 42306 41064
rect 44192 41052 44220 41083
rect 45002 41080 45008 41132
rect 45060 41120 45066 41132
rect 45097 41123 45155 41129
rect 45097 41120 45109 41123
rect 45060 41092 45109 41120
rect 45060 41080 45066 41092
rect 45097 41089 45109 41092
rect 45143 41120 45155 41123
rect 45738 41120 45744 41132
rect 45143 41092 45744 41120
rect 45143 41089 45155 41092
rect 45097 41083 45155 41089
rect 45738 41080 45744 41092
rect 45796 41080 45802 41132
rect 46014 41080 46020 41132
rect 46072 41120 46078 41132
rect 46290 41120 46296 41132
rect 46072 41092 46296 41120
rect 46072 41080 46078 41092
rect 46290 41080 46296 41092
rect 46348 41120 46354 41132
rect 50890 41120 50896 41132
rect 46348 41092 50896 41120
rect 46348 41080 46354 41092
rect 50890 41080 50896 41092
rect 50948 41080 50954 41132
rect 51046 41120 51074 41228
rect 51350 41216 51356 41268
rect 51408 41216 51414 41268
rect 53098 41216 53104 41268
rect 53156 41256 53162 41268
rect 54018 41256 54024 41268
rect 53156 41228 54024 41256
rect 53156 41216 53162 41228
rect 54018 41216 54024 41228
rect 54076 41216 54082 41268
rect 56502 41216 56508 41268
rect 56560 41216 56566 41268
rect 58066 41148 58072 41200
rect 58124 41188 58130 41200
rect 66438 41188 66444 41200
rect 58124 41160 66444 41188
rect 58124 41148 58130 41160
rect 66438 41148 66444 41160
rect 66496 41148 66502 41200
rect 51046 41092 51212 41120
rect 44266 41052 44272 41064
rect 44192 41024 44272 41052
rect 44266 41012 44272 41024
rect 44324 41052 44330 41064
rect 44821 41055 44879 41061
rect 44821 41052 44833 41055
rect 44324 41024 44833 41052
rect 44324 41012 44330 41024
rect 44821 41021 44833 41024
rect 44867 41052 44879 41055
rect 46753 41055 46811 41061
rect 46753 41052 46765 41055
rect 44867 41024 46765 41052
rect 44867 41021 44879 41024
rect 44821 41015 44879 41021
rect 46753 41021 46765 41024
rect 46799 41021 46811 41055
rect 46753 41015 46811 41021
rect 46934 41012 46940 41064
rect 46992 41012 46998 41064
rect 48314 41012 48320 41064
rect 48372 41012 48378 41064
rect 49602 41012 49608 41064
rect 49660 41012 49666 41064
rect 51184 41052 51212 41092
rect 52638 41080 52644 41132
rect 52696 41120 52702 41132
rect 53837 41123 53895 41129
rect 53837 41120 53849 41123
rect 52696 41092 53849 41120
rect 52696 41080 52702 41092
rect 53837 41089 53849 41092
rect 53883 41089 53895 41123
rect 53837 41083 53895 41089
rect 53926 41080 53932 41132
rect 53984 41120 53990 41132
rect 54110 41120 54116 41132
rect 53984 41092 54116 41120
rect 53984 41080 53990 41092
rect 54110 41080 54116 41092
rect 54168 41080 54174 41132
rect 64874 41120 64880 41132
rect 54404 41092 64880 41120
rect 51445 41055 51503 41061
rect 51445 41052 51457 41055
rect 51184 41024 51457 41052
rect 51445 41021 51457 41024
rect 51491 41052 51503 41055
rect 54404 41052 54432 41092
rect 64874 41080 64880 41092
rect 64932 41080 64938 41132
rect 51491 41024 54432 41052
rect 51491 41021 51503 41024
rect 51445 41015 51503 41021
rect 54754 41012 54760 41064
rect 54812 41012 54818 41064
rect 56686 41012 56692 41064
rect 56744 41052 56750 41064
rect 56965 41055 57023 41061
rect 56965 41052 56977 41055
rect 56744 41024 56977 41052
rect 56744 41012 56750 41024
rect 56965 41021 56977 41024
rect 57011 41052 57023 41055
rect 57149 41055 57207 41061
rect 57149 41052 57161 41055
rect 57011 41024 57161 41052
rect 57011 41021 57023 41024
rect 56965 41015 57023 41021
rect 57149 41021 57161 41024
rect 57195 41021 57207 41055
rect 57149 41015 57207 41021
rect 57241 41055 57299 41061
rect 57241 41021 57253 41055
rect 57287 41021 57299 41055
rect 57241 41015 57299 41021
rect 33778 40984 33784 40996
rect 33612 40956 33784 40984
rect 33505 40947 33563 40953
rect 33778 40944 33784 40956
rect 33836 40944 33842 40996
rect 35161 40987 35219 40993
rect 35161 40953 35173 40987
rect 35207 40953 35219 40987
rect 35161 40947 35219 40953
rect 38488 40956 40448 40984
rect 22186 40916 22192 40928
rect 20220 40888 22192 40916
rect 20220 40876 20226 40888
rect 22186 40876 22192 40888
rect 22244 40876 22250 40928
rect 23750 40876 23756 40928
rect 23808 40916 23814 40928
rect 23845 40919 23903 40925
rect 23845 40916 23857 40919
rect 23808 40888 23857 40916
rect 23808 40876 23814 40888
rect 23845 40885 23857 40888
rect 23891 40885 23903 40919
rect 23845 40879 23903 40885
rect 24305 40919 24363 40925
rect 24305 40885 24317 40919
rect 24351 40916 24363 40919
rect 25130 40916 25136 40928
rect 24351 40888 25136 40916
rect 24351 40885 24363 40888
rect 24305 40879 24363 40885
rect 25130 40876 25136 40888
rect 25188 40876 25194 40928
rect 26145 40919 26203 40925
rect 26145 40885 26157 40919
rect 26191 40916 26203 40919
rect 26234 40916 26240 40928
rect 26191 40888 26240 40916
rect 26191 40885 26203 40888
rect 26145 40879 26203 40885
rect 26234 40876 26240 40888
rect 26292 40876 26298 40928
rect 29454 40876 29460 40928
rect 29512 40876 29518 40928
rect 29825 40919 29883 40925
rect 29825 40885 29837 40919
rect 29871 40916 29883 40919
rect 29914 40916 29920 40928
rect 29871 40888 29920 40916
rect 29871 40885 29883 40888
rect 29825 40879 29883 40885
rect 29914 40876 29920 40888
rect 29972 40876 29978 40928
rect 30006 40876 30012 40928
rect 30064 40916 30070 40928
rect 30466 40916 30472 40928
rect 30064 40888 30472 40916
rect 30064 40876 30070 40888
rect 30466 40876 30472 40888
rect 30524 40876 30530 40928
rect 31018 40876 31024 40928
rect 31076 40916 31082 40928
rect 31297 40919 31355 40925
rect 31297 40916 31309 40919
rect 31076 40888 31309 40916
rect 31076 40876 31082 40888
rect 31297 40885 31309 40888
rect 31343 40885 31355 40919
rect 31297 40879 31355 40885
rect 31386 40876 31392 40928
rect 31444 40916 31450 40928
rect 32950 40916 32956 40928
rect 31444 40888 32956 40916
rect 31444 40876 31450 40888
rect 32950 40876 32956 40888
rect 33008 40876 33014 40928
rect 33042 40876 33048 40928
rect 33100 40916 33106 40928
rect 33137 40919 33195 40925
rect 33137 40916 33149 40919
rect 33100 40888 33149 40916
rect 33100 40876 33106 40888
rect 33137 40885 33149 40888
rect 33183 40885 33195 40919
rect 33137 40879 33195 40885
rect 33594 40876 33600 40928
rect 33652 40876 33658 40928
rect 33962 40876 33968 40928
rect 34020 40916 34026 40928
rect 34149 40919 34207 40925
rect 34149 40916 34161 40919
rect 34020 40888 34161 40916
rect 34020 40876 34026 40888
rect 34149 40885 34161 40888
rect 34195 40885 34207 40919
rect 35176 40916 35204 40947
rect 35802 40916 35808 40928
rect 35176 40888 35808 40916
rect 34149 40879 34207 40885
rect 35802 40876 35808 40888
rect 35860 40876 35866 40928
rect 36998 40876 37004 40928
rect 37056 40916 37062 40928
rect 37277 40919 37335 40925
rect 37277 40916 37289 40919
rect 37056 40888 37289 40916
rect 37056 40876 37062 40888
rect 37277 40885 37289 40888
rect 37323 40885 37335 40919
rect 37277 40879 37335 40885
rect 37645 40919 37703 40925
rect 37645 40885 37657 40919
rect 37691 40916 37703 40919
rect 37826 40916 37832 40928
rect 37691 40888 37832 40916
rect 37691 40885 37703 40888
rect 37645 40879 37703 40885
rect 37826 40876 37832 40888
rect 37884 40876 37890 40928
rect 38102 40876 38108 40928
rect 38160 40876 38166 40928
rect 38488 40925 38516 40956
rect 38473 40919 38531 40925
rect 38473 40885 38485 40919
rect 38519 40885 38531 40919
rect 38473 40879 38531 40885
rect 38565 40919 38623 40925
rect 38565 40885 38577 40919
rect 38611 40916 38623 40919
rect 39206 40916 39212 40928
rect 38611 40888 39212 40916
rect 38611 40885 38623 40888
rect 38565 40879 38623 40885
rect 39206 40876 39212 40888
rect 39264 40876 39270 40928
rect 39301 40919 39359 40925
rect 39301 40885 39313 40919
rect 39347 40916 39359 40919
rect 39482 40916 39488 40928
rect 39347 40888 39488 40916
rect 39347 40885 39359 40888
rect 39301 40879 39359 40885
rect 39482 40876 39488 40888
rect 39540 40876 39546 40928
rect 39666 40876 39672 40928
rect 39724 40876 39730 40928
rect 40420 40916 40448 40956
rect 40494 40944 40500 40996
rect 40552 40944 40558 40996
rect 42610 40944 42616 40996
rect 42668 40984 42674 40996
rect 42705 40987 42763 40993
rect 42705 40984 42717 40987
rect 42668 40956 42717 40984
rect 42668 40944 42674 40956
rect 42705 40953 42717 40956
rect 42751 40953 42763 40987
rect 42705 40947 42763 40953
rect 42794 40944 42800 40996
rect 42852 40984 42858 40996
rect 43162 40984 43168 40996
rect 42852 40956 43168 40984
rect 42852 40944 42858 40956
rect 43162 40944 43168 40956
rect 43220 40944 43226 40996
rect 44913 40987 44971 40993
rect 44913 40953 44925 40987
rect 44959 40984 44971 40987
rect 46014 40984 46020 40996
rect 44959 40956 46020 40984
rect 44959 40953 44971 40956
rect 44913 40947 44971 40953
rect 46014 40944 46020 40956
rect 46072 40944 46078 40996
rect 47210 40944 47216 40996
rect 47268 40944 47274 40996
rect 49786 40944 49792 40996
rect 49844 40984 49850 40996
rect 49881 40987 49939 40993
rect 49881 40984 49893 40987
rect 49844 40956 49893 40984
rect 49844 40944 49850 40956
rect 49881 40953 49893 40956
rect 49927 40953 49939 40987
rect 50338 40984 50344 40996
rect 49881 40947 49939 40953
rect 49988 40956 50344 40984
rect 41046 40916 41052 40928
rect 40420 40888 41052 40916
rect 41046 40876 41052 40888
rect 41104 40876 41110 40928
rect 45094 40876 45100 40928
rect 45152 40916 45158 40928
rect 45373 40919 45431 40925
rect 45373 40916 45385 40919
rect 45152 40888 45385 40916
rect 45152 40876 45158 40888
rect 45373 40885 45385 40888
rect 45419 40885 45431 40919
rect 45373 40879 45431 40885
rect 45738 40876 45744 40928
rect 45796 40876 45802 40928
rect 45830 40876 45836 40928
rect 45888 40876 45894 40928
rect 48222 40876 48228 40928
rect 48280 40916 48286 40928
rect 48682 40916 48688 40928
rect 48280 40888 48688 40916
rect 48280 40876 48286 40888
rect 48682 40876 48688 40888
rect 48740 40876 48746 40928
rect 48958 40876 48964 40928
rect 49016 40916 49022 40928
rect 49988 40916 50016 40956
rect 50338 40944 50344 40956
rect 50396 40944 50402 40996
rect 52178 40944 52184 40996
rect 52236 40984 52242 40996
rect 53193 40987 53251 40993
rect 53193 40984 53205 40987
rect 52236 40956 53205 40984
rect 52236 40944 52242 40956
rect 53193 40953 53205 40956
rect 53239 40984 53251 40987
rect 54772 40984 54800 41012
rect 53239 40956 54800 40984
rect 53239 40953 53251 40956
rect 53193 40947 53251 40953
rect 55030 40944 55036 40996
rect 55088 40944 55094 40996
rect 55122 40944 55128 40996
rect 55180 40984 55186 40996
rect 55180 40956 55522 40984
rect 55180 40944 55186 40956
rect 56594 40944 56600 40996
rect 56652 40944 56658 40996
rect 57256 40984 57284 41015
rect 57422 41012 57428 41064
rect 57480 41012 57486 41064
rect 57164 40956 57284 40984
rect 49016 40888 50016 40916
rect 53285 40919 53343 40925
rect 49016 40876 49022 40888
rect 53285 40885 53297 40919
rect 53331 40916 53343 40919
rect 53466 40916 53472 40928
rect 53331 40888 53472 40916
rect 53331 40885 53343 40888
rect 53285 40879 53343 40885
rect 53466 40876 53472 40888
rect 53524 40876 53530 40928
rect 53650 40876 53656 40928
rect 53708 40876 53714 40928
rect 53745 40919 53803 40925
rect 53745 40885 53757 40919
rect 53791 40916 53803 40919
rect 53926 40916 53932 40928
rect 53791 40888 53932 40916
rect 53791 40885 53803 40888
rect 53745 40879 53803 40885
rect 53926 40876 53932 40888
rect 53984 40876 53990 40928
rect 54110 40876 54116 40928
rect 54168 40916 54174 40928
rect 54662 40916 54668 40928
rect 54168 40888 54668 40916
rect 54168 40876 54174 40888
rect 54662 40876 54668 40888
rect 54720 40916 54726 40928
rect 57164 40916 57192 40956
rect 54720 40888 57192 40916
rect 54720 40876 54726 40888
rect 552 40826 66424 40848
rect 552 40774 2918 40826
rect 2970 40774 2982 40826
rect 3034 40774 3046 40826
rect 3098 40774 3110 40826
rect 3162 40774 3174 40826
rect 3226 40774 50918 40826
rect 50970 40774 50982 40826
rect 51034 40774 51046 40826
rect 51098 40774 51110 40826
rect 51162 40774 51174 40826
rect 51226 40774 66424 40826
rect 552 40752 66424 40774
rect 7929 40715 7987 40721
rect 7929 40681 7941 40715
rect 7975 40712 7987 40715
rect 8018 40712 8024 40724
rect 7975 40684 8024 40712
rect 7975 40681 7987 40684
rect 7929 40675 7987 40681
rect 8018 40672 8024 40684
rect 8076 40672 8082 40724
rect 8297 40715 8355 40721
rect 8297 40681 8309 40715
rect 8343 40712 8355 40715
rect 8938 40712 8944 40724
rect 8343 40684 8944 40712
rect 8343 40681 8355 40684
rect 8297 40675 8355 40681
rect 8938 40672 8944 40684
rect 8996 40672 9002 40724
rect 11330 40672 11336 40724
rect 11388 40712 11394 40724
rect 13998 40712 14004 40724
rect 11388 40684 14004 40712
rect 11388 40672 11394 40684
rect 13998 40672 14004 40684
rect 14056 40672 14062 40724
rect 15194 40672 15200 40724
rect 15252 40672 15258 40724
rect 15470 40672 15476 40724
rect 15528 40712 15534 40724
rect 15565 40715 15623 40721
rect 15565 40712 15577 40715
rect 15528 40684 15577 40712
rect 15528 40672 15534 40684
rect 15565 40681 15577 40684
rect 15611 40681 15623 40715
rect 15565 40675 15623 40681
rect 15657 40715 15715 40721
rect 15657 40681 15669 40715
rect 15703 40712 15715 40715
rect 17402 40712 17408 40724
rect 15703 40684 17408 40712
rect 15703 40681 15715 40684
rect 15657 40675 15715 40681
rect 17402 40672 17408 40684
rect 17460 40672 17466 40724
rect 17770 40672 17776 40724
rect 17828 40712 17834 40724
rect 17828 40684 21956 40712
rect 17828 40672 17834 40684
rect 9030 40604 9036 40656
rect 9088 40604 9094 40656
rect 10318 40644 10324 40656
rect 10258 40616 10324 40644
rect 10318 40604 10324 40616
rect 10376 40644 10382 40656
rect 10962 40644 10968 40656
rect 10376 40616 10968 40644
rect 10376 40604 10382 40616
rect 10962 40604 10968 40616
rect 11020 40604 11026 40656
rect 12434 40604 12440 40656
rect 12492 40604 12498 40656
rect 12526 40604 12532 40656
rect 12584 40644 12590 40656
rect 12584 40616 12926 40644
rect 12584 40604 12590 40616
rect 15010 40604 15016 40656
rect 15068 40644 15074 40656
rect 15068 40616 16160 40644
rect 15068 40604 15074 40616
rect 8294 40536 8300 40588
rect 8352 40576 8358 40588
rect 8352 40548 8616 40576
rect 8352 40536 8358 40548
rect 8588 40520 8616 40548
rect 10778 40536 10784 40588
rect 10836 40576 10842 40588
rect 11425 40579 11483 40585
rect 11425 40576 11437 40579
rect 10836 40548 11437 40576
rect 10836 40536 10842 40548
rect 11425 40545 11437 40548
rect 11471 40576 11483 40579
rect 11698 40576 11704 40588
rect 11471 40548 11704 40576
rect 11471 40545 11483 40548
rect 11425 40539 11483 40545
rect 11698 40536 11704 40548
rect 11756 40536 11762 40588
rect 14550 40536 14556 40588
rect 14608 40536 14614 40588
rect 15838 40576 15844 40588
rect 15212 40548 15844 40576
rect 8389 40511 8447 40517
rect 8389 40477 8401 40511
rect 8435 40477 8447 40511
rect 8389 40471 8447 40477
rect 8404 40440 8432 40471
rect 8570 40468 8576 40520
rect 8628 40468 8634 40520
rect 8754 40468 8760 40520
rect 8812 40468 8818 40520
rect 10410 40508 10416 40520
rect 8864 40480 10416 40508
rect 8864 40440 8892 40480
rect 10410 40468 10416 40480
rect 10468 40468 10474 40520
rect 11238 40468 11244 40520
rect 11296 40508 11302 40520
rect 11517 40511 11575 40517
rect 11517 40508 11529 40511
rect 11296 40480 11529 40508
rect 11296 40468 11302 40480
rect 11517 40477 11529 40480
rect 11563 40508 11575 40511
rect 12066 40508 12072 40520
rect 11563 40480 12072 40508
rect 11563 40477 11575 40480
rect 11517 40471 11575 40477
rect 12066 40468 12072 40480
rect 12124 40468 12130 40520
rect 12161 40511 12219 40517
rect 12161 40477 12173 40511
rect 12207 40508 12219 40511
rect 13814 40508 13820 40520
rect 12207 40480 13820 40508
rect 12207 40477 12219 40480
rect 12161 40471 12219 40477
rect 8404 40412 8892 40440
rect 10686 40400 10692 40452
rect 10744 40440 10750 40452
rect 12176 40440 12204 40471
rect 13814 40468 13820 40480
rect 13872 40468 13878 40520
rect 13906 40468 13912 40520
rect 13964 40508 13970 40520
rect 14185 40511 14243 40517
rect 14185 40508 14197 40511
rect 13964 40480 14197 40508
rect 13964 40468 13970 40480
rect 14185 40477 14197 40480
rect 14231 40508 14243 40511
rect 15212 40508 15240 40548
rect 15838 40536 15844 40548
rect 15896 40536 15902 40588
rect 16132 40585 16160 40616
rect 16850 40604 16856 40656
rect 16908 40604 16914 40656
rect 21818 40644 21824 40656
rect 21560 40616 21824 40644
rect 16117 40579 16175 40585
rect 16117 40545 16129 40579
rect 16163 40545 16175 40579
rect 16117 40539 16175 40545
rect 18049 40579 18107 40585
rect 18049 40545 18061 40579
rect 18095 40576 18107 40579
rect 18506 40576 18512 40588
rect 18095 40548 18512 40576
rect 18095 40545 18107 40548
rect 18049 40539 18107 40545
rect 18506 40536 18512 40548
rect 18564 40536 18570 40588
rect 19242 40536 19248 40588
rect 19300 40576 19306 40588
rect 21560 40576 21588 40616
rect 21818 40604 21824 40616
rect 21876 40604 21882 40656
rect 21928 40644 21956 40684
rect 22002 40672 22008 40724
rect 22060 40672 22066 40724
rect 22925 40715 22983 40721
rect 22925 40681 22937 40715
rect 22971 40712 22983 40715
rect 23014 40712 23020 40724
rect 22971 40684 23020 40712
rect 22971 40681 22983 40684
rect 22925 40675 22983 40681
rect 23014 40672 23020 40684
rect 23072 40672 23078 40724
rect 26234 40712 26240 40724
rect 23492 40684 26240 40712
rect 21928 40616 23060 40644
rect 19300 40548 19642 40576
rect 21468 40548 21588 40576
rect 21637 40579 21695 40585
rect 19300 40536 19306 40548
rect 21468 40520 21496 40548
rect 21637 40545 21649 40579
rect 21683 40576 21695 40579
rect 22646 40576 22652 40588
rect 21683 40548 22652 40576
rect 21683 40545 21695 40548
rect 21637 40539 21695 40545
rect 22646 40536 22652 40548
rect 22704 40536 22710 40588
rect 14231 40480 15240 40508
rect 14231 40477 14243 40480
rect 14185 40471 14243 40477
rect 15286 40468 15292 40520
rect 15344 40508 15350 40520
rect 15654 40508 15660 40520
rect 15344 40480 15660 40508
rect 15344 40468 15350 40480
rect 15654 40468 15660 40480
rect 15712 40508 15718 40520
rect 15749 40511 15807 40517
rect 15749 40508 15761 40511
rect 15712 40480 15761 40508
rect 15712 40468 15718 40480
rect 15749 40477 15761 40480
rect 15795 40477 15807 40511
rect 15749 40471 15807 40477
rect 15930 40468 15936 40520
rect 15988 40508 15994 40520
rect 16393 40511 16451 40517
rect 16393 40508 16405 40511
rect 15988 40480 16405 40508
rect 15988 40468 15994 40480
rect 16393 40477 16405 40480
rect 16439 40477 16451 40511
rect 16393 40471 16451 40477
rect 16482 40468 16488 40520
rect 16540 40508 16546 40520
rect 18601 40511 18659 40517
rect 18601 40508 18613 40511
rect 16540 40480 18613 40508
rect 16540 40468 16546 40480
rect 18601 40477 18613 40480
rect 18647 40477 18659 40511
rect 18601 40471 18659 40477
rect 18782 40468 18788 40520
rect 18840 40468 18846 40520
rect 20714 40468 20720 40520
rect 20772 40468 20778 40520
rect 20993 40511 21051 40517
rect 20993 40477 21005 40511
rect 21039 40477 21051 40511
rect 20993 40471 21051 40477
rect 10744 40412 12204 40440
rect 10744 40400 10750 40412
rect 17402 40400 17408 40452
rect 17460 40440 17466 40452
rect 18141 40443 18199 40449
rect 18141 40440 18153 40443
rect 17460 40412 18153 40440
rect 17460 40400 17466 40412
rect 18141 40409 18153 40412
rect 18187 40409 18199 40443
rect 18141 40403 18199 40409
rect 18322 40400 18328 40452
rect 18380 40440 18386 40452
rect 21008 40440 21036 40471
rect 21450 40468 21456 40520
rect 21508 40468 21514 40520
rect 21542 40468 21548 40520
rect 21600 40468 21606 40520
rect 21726 40468 21732 40520
rect 21784 40508 21790 40520
rect 22097 40511 22155 40517
rect 22097 40508 22109 40511
rect 21784 40480 22109 40508
rect 21784 40468 21790 40480
rect 22097 40477 22109 40480
rect 22143 40477 22155 40511
rect 23032 40508 23060 40616
rect 23198 40604 23204 40656
rect 23256 40604 23262 40656
rect 23492 40585 23520 40684
rect 26234 40672 26240 40684
rect 26292 40672 26298 40724
rect 26510 40672 26516 40724
rect 26568 40712 26574 40724
rect 26568 40684 27384 40712
rect 26568 40672 26574 40684
rect 23750 40604 23756 40656
rect 23808 40604 23814 40656
rect 25685 40647 25743 40653
rect 25685 40613 25697 40647
rect 25731 40644 25743 40647
rect 27246 40644 27252 40656
rect 25731 40616 27252 40644
rect 25731 40613 25743 40616
rect 25685 40607 25743 40613
rect 23477 40579 23535 40585
rect 23477 40545 23489 40579
rect 23523 40545 23535 40579
rect 23477 40539 23535 40545
rect 24762 40508 24768 40520
rect 23032 40480 24768 40508
rect 22097 40471 22155 40477
rect 24762 40468 24768 40480
rect 24820 40468 24826 40520
rect 24872 40508 24900 40562
rect 24946 40508 24952 40520
rect 24872 40480 24952 40508
rect 24946 40468 24952 40480
rect 25004 40468 25010 40520
rect 25225 40511 25283 40517
rect 25225 40477 25237 40511
rect 25271 40508 25283 40511
rect 25700 40508 25728 40607
rect 27246 40604 27252 40616
rect 27304 40604 27310 40656
rect 27356 40585 27384 40684
rect 27430 40672 27436 40724
rect 27488 40712 27494 40724
rect 28258 40712 28264 40724
rect 27488 40684 28264 40712
rect 27488 40672 27494 40684
rect 28258 40672 28264 40684
rect 28316 40672 28322 40724
rect 29457 40715 29515 40721
rect 29457 40681 29469 40715
rect 29503 40681 29515 40715
rect 29457 40675 29515 40681
rect 25777 40579 25835 40585
rect 25777 40545 25789 40579
rect 25823 40576 25835 40579
rect 26421 40579 26479 40585
rect 26421 40576 26433 40579
rect 25823 40548 26433 40576
rect 25823 40545 25835 40548
rect 25777 40539 25835 40545
rect 26421 40545 26433 40548
rect 26467 40545 26479 40579
rect 26421 40539 26479 40545
rect 27341 40579 27399 40585
rect 27341 40545 27353 40579
rect 27387 40576 27399 40579
rect 27617 40579 27675 40585
rect 27617 40576 27629 40579
rect 27387 40548 27629 40576
rect 27387 40545 27399 40548
rect 27341 40539 27399 40545
rect 27617 40545 27629 40548
rect 27663 40545 27675 40579
rect 27617 40539 27675 40545
rect 28994 40536 29000 40588
rect 29052 40536 29058 40588
rect 25271 40480 25728 40508
rect 25961 40511 26019 40517
rect 25271 40477 25283 40480
rect 25225 40471 25283 40477
rect 25961 40477 25973 40511
rect 26007 40508 26019 40511
rect 26050 40508 26056 40520
rect 26007 40480 26056 40508
rect 26007 40477 26019 40480
rect 25961 40471 26019 40477
rect 26050 40468 26056 40480
rect 26108 40468 26114 40520
rect 27062 40468 27068 40520
rect 27120 40468 27126 40520
rect 27893 40511 27951 40517
rect 27893 40477 27905 40511
rect 27939 40508 27951 40511
rect 29472 40508 29500 40675
rect 29914 40672 29920 40724
rect 29972 40672 29978 40724
rect 31018 40672 31024 40724
rect 31076 40672 31082 40724
rect 32214 40672 32220 40724
rect 32272 40672 32278 40724
rect 32766 40672 32772 40724
rect 32824 40712 32830 40724
rect 33505 40715 33563 40721
rect 32824 40684 33364 40712
rect 32824 40672 32830 40684
rect 32232 40644 32260 40672
rect 31772 40616 32260 40644
rect 33336 40644 33364 40684
rect 33505 40681 33517 40715
rect 33551 40712 33563 40715
rect 33686 40712 33692 40724
rect 33551 40684 33692 40712
rect 33551 40681 33563 40684
rect 33505 40675 33563 40681
rect 33686 40672 33692 40684
rect 33744 40672 33750 40724
rect 33962 40672 33968 40724
rect 34020 40672 34026 40724
rect 36170 40712 36176 40724
rect 34072 40684 36176 40712
rect 34072 40644 34100 40684
rect 36170 40672 36176 40684
rect 36228 40672 36234 40724
rect 36722 40672 36728 40724
rect 36780 40712 36786 40724
rect 37185 40715 37243 40721
rect 37185 40712 37197 40715
rect 36780 40684 37197 40712
rect 36780 40672 36786 40684
rect 37185 40681 37197 40684
rect 37231 40712 37243 40715
rect 37918 40712 37924 40724
rect 37231 40684 37924 40712
rect 37231 40681 37243 40684
rect 37185 40675 37243 40681
rect 37918 40672 37924 40684
rect 37976 40672 37982 40724
rect 40494 40712 40500 40724
rect 39224 40684 40500 40712
rect 33336 40616 34100 40644
rect 31772 40588 31800 40616
rect 34790 40604 34796 40656
rect 34848 40604 34854 40656
rect 36538 40604 36544 40656
rect 36596 40644 36602 40656
rect 38470 40644 38476 40656
rect 36596 40616 38476 40644
rect 36596 40604 36602 40616
rect 38470 40604 38476 40616
rect 38528 40604 38534 40656
rect 29822 40536 29828 40588
rect 29880 40536 29886 40588
rect 30834 40576 30840 40588
rect 30116 40548 30840 40576
rect 30116 40517 30144 40548
rect 30834 40536 30840 40548
rect 30892 40576 30898 40588
rect 31662 40576 31668 40588
rect 30892 40548 31668 40576
rect 30892 40536 30898 40548
rect 31662 40536 31668 40548
rect 31720 40536 31726 40588
rect 31754 40536 31760 40588
rect 31812 40536 31818 40588
rect 33134 40536 33140 40588
rect 33192 40576 33198 40588
rect 36078 40576 36084 40588
rect 33192 40548 36084 40576
rect 33192 40536 33198 40548
rect 36078 40536 36084 40548
rect 36136 40536 36142 40588
rect 39224 40585 39252 40684
rect 40494 40672 40500 40684
rect 40552 40672 40558 40724
rect 41046 40672 41052 40724
rect 41104 40672 41110 40724
rect 41506 40672 41512 40724
rect 41564 40712 41570 40724
rect 42058 40712 42064 40724
rect 41564 40684 42064 40712
rect 41564 40672 41570 40684
rect 42058 40672 42064 40684
rect 42116 40672 42122 40724
rect 42242 40672 42248 40724
rect 42300 40712 42306 40724
rect 65058 40712 65064 40724
rect 42300 40684 65064 40712
rect 42300 40672 42306 40684
rect 39482 40604 39488 40656
rect 39540 40604 39546 40656
rect 40954 40644 40960 40656
rect 40710 40616 40960 40644
rect 40954 40604 40960 40616
rect 41012 40604 41018 40656
rect 42613 40647 42671 40653
rect 42613 40613 42625 40647
rect 42659 40644 42671 40647
rect 42886 40644 42892 40656
rect 42659 40616 42892 40644
rect 42659 40613 42671 40616
rect 42613 40607 42671 40613
rect 42886 40604 42892 40616
rect 42944 40604 42950 40656
rect 43162 40604 43168 40656
rect 43220 40604 43226 40656
rect 45094 40604 45100 40656
rect 45152 40604 45158 40656
rect 46474 40644 46480 40656
rect 46322 40616 46480 40644
rect 46474 40604 46480 40616
rect 46532 40604 46538 40656
rect 47762 40604 47768 40656
rect 47820 40604 47826 40656
rect 47946 40604 47952 40656
rect 48004 40644 48010 40656
rect 49694 40644 49700 40656
rect 48004 40616 49700 40644
rect 48004 40604 48010 40616
rect 39209 40579 39267 40585
rect 39209 40545 39221 40579
rect 39255 40545 39267 40579
rect 39209 40539 39267 40545
rect 41966 40536 41972 40588
rect 42024 40576 42030 40588
rect 42242 40576 42248 40588
rect 42024 40548 42248 40576
rect 42024 40536 42030 40548
rect 42242 40536 42248 40548
rect 42300 40536 42306 40588
rect 47854 40536 47860 40588
rect 47912 40536 47918 40588
rect 27939 40480 29500 40508
rect 30101 40511 30159 40517
rect 27939 40477 27951 40480
rect 27893 40471 27951 40477
rect 30101 40477 30113 40511
rect 30147 40477 30159 40511
rect 30101 40471 30159 40477
rect 31110 40468 31116 40520
rect 31168 40468 31174 40520
rect 31294 40468 31300 40520
rect 31352 40468 31358 40520
rect 32033 40511 32091 40517
rect 32033 40477 32045 40511
rect 32079 40508 32091 40511
rect 32079 40480 33640 40508
rect 32079 40477 32091 40480
rect 32033 40471 32091 40477
rect 22186 40440 22192 40452
rect 18380 40412 19472 40440
rect 21008 40412 22192 40440
rect 18380 40400 18386 40412
rect 7742 40332 7748 40384
rect 7800 40372 7806 40384
rect 10965 40375 11023 40381
rect 10965 40372 10977 40375
rect 7800 40344 10977 40372
rect 7800 40332 7806 40344
rect 10965 40341 10977 40344
rect 11011 40341 11023 40375
rect 10965 40335 11023 40341
rect 15105 40375 15163 40381
rect 15105 40341 15117 40375
rect 15151 40372 15163 40375
rect 15562 40372 15568 40384
rect 15151 40344 15568 40372
rect 15151 40341 15163 40344
rect 15105 40335 15163 40341
rect 15562 40332 15568 40344
rect 15620 40332 15626 40384
rect 15746 40332 15752 40384
rect 15804 40372 15810 40384
rect 16850 40372 16856 40384
rect 15804 40344 16856 40372
rect 15804 40332 15810 40344
rect 16850 40332 16856 40344
rect 16908 40372 16914 40384
rect 17678 40372 17684 40384
rect 16908 40344 17684 40372
rect 16908 40332 16914 40344
rect 17678 40332 17684 40344
rect 17736 40332 17742 40384
rect 17862 40332 17868 40384
rect 17920 40332 17926 40384
rect 19245 40375 19303 40381
rect 19245 40341 19257 40375
rect 19291 40372 19303 40375
rect 19334 40372 19340 40384
rect 19291 40344 19340 40372
rect 19291 40341 19303 40344
rect 19245 40335 19303 40341
rect 19334 40332 19340 40344
rect 19392 40332 19398 40384
rect 19444 40372 19472 40412
rect 22186 40400 22192 40412
rect 22244 40400 22250 40452
rect 23014 40440 23020 40452
rect 22480 40412 23020 40440
rect 21450 40372 21456 40384
rect 19444 40344 21456 40372
rect 21450 40332 21456 40344
rect 21508 40332 21514 40384
rect 21634 40332 21640 40384
rect 21692 40372 21698 40384
rect 22002 40372 22008 40384
rect 21692 40344 22008 40372
rect 21692 40332 21698 40344
rect 22002 40332 22008 40344
rect 22060 40372 22066 40384
rect 22480 40372 22508 40412
rect 23014 40400 23020 40412
rect 23072 40400 23078 40452
rect 25038 40400 25044 40452
rect 25096 40440 25102 40452
rect 27522 40440 27528 40452
rect 25096 40412 27528 40440
rect 25096 40400 25102 40412
rect 27522 40400 27528 40412
rect 27580 40400 27586 40452
rect 33502 40440 33508 40452
rect 28920 40412 31754 40440
rect 22060 40344 22508 40372
rect 22060 40332 22066 40344
rect 22738 40332 22744 40384
rect 22796 40332 22802 40384
rect 25314 40332 25320 40384
rect 25372 40332 25378 40384
rect 26602 40332 26608 40384
rect 26660 40372 26666 40384
rect 28920 40372 28948 40412
rect 26660 40344 28948 40372
rect 26660 40332 26666 40344
rect 29362 40332 29368 40384
rect 29420 40372 29426 40384
rect 30558 40372 30564 40384
rect 29420 40344 30564 40372
rect 29420 40332 29426 40344
rect 30558 40332 30564 40344
rect 30616 40332 30622 40384
rect 30650 40332 30656 40384
rect 30708 40332 30714 40384
rect 31726 40372 31754 40412
rect 33152 40412 33508 40440
rect 33152 40372 33180 40412
rect 33502 40400 33508 40412
rect 33560 40400 33566 40452
rect 33612 40449 33640 40480
rect 34054 40468 34060 40520
rect 34112 40468 34118 40520
rect 34146 40468 34152 40520
rect 34204 40468 34210 40520
rect 39850 40468 39856 40520
rect 39908 40508 39914 40520
rect 41601 40511 41659 40517
rect 41601 40508 41613 40511
rect 39908 40480 41613 40508
rect 39908 40468 39914 40480
rect 41601 40477 41613 40480
rect 41647 40477 41659 40511
rect 41601 40471 41659 40477
rect 41874 40468 41880 40520
rect 41932 40508 41938 40520
rect 42337 40511 42395 40517
rect 42337 40508 42349 40511
rect 41932 40480 42349 40508
rect 41932 40468 41938 40480
rect 42337 40477 42349 40480
rect 42383 40477 42395 40511
rect 44818 40508 44824 40520
rect 42337 40471 42395 40477
rect 42444 40480 44824 40508
rect 33597 40443 33655 40449
rect 33597 40409 33609 40443
rect 33643 40409 33655 40443
rect 33597 40403 33655 40409
rect 34882 40400 34888 40452
rect 34940 40440 34946 40452
rect 36081 40443 36139 40449
rect 36081 40440 36093 40443
rect 34940 40412 36093 40440
rect 34940 40400 34946 40412
rect 36081 40409 36093 40412
rect 36127 40440 36139 40443
rect 37366 40440 37372 40452
rect 36127 40412 37372 40440
rect 36127 40409 36139 40412
rect 36081 40403 36139 40409
rect 37366 40400 37372 40412
rect 37424 40440 37430 40452
rect 37734 40440 37740 40452
rect 37424 40412 37740 40440
rect 37424 40400 37430 40412
rect 37734 40400 37740 40412
rect 37792 40400 37798 40452
rect 41690 40400 41696 40452
rect 41748 40440 41754 40452
rect 42444 40440 42472 40480
rect 44818 40468 44824 40480
rect 44876 40468 44882 40520
rect 48056 40517 48084 40616
rect 49694 40604 49700 40616
rect 49752 40604 49758 40656
rect 50264 40653 50292 40684
rect 65058 40672 65064 40684
rect 65116 40672 65122 40724
rect 50249 40647 50307 40653
rect 50249 40613 50261 40647
rect 50295 40613 50307 40647
rect 50249 40607 50307 40613
rect 52454 40604 52460 40656
rect 52512 40604 52518 40656
rect 53098 40604 53104 40656
rect 53156 40604 53162 40656
rect 54018 40604 54024 40656
rect 54076 40644 54082 40656
rect 55122 40644 55128 40656
rect 54076 40616 55128 40644
rect 54076 40604 54082 40616
rect 55122 40604 55128 40616
rect 55180 40644 55186 40656
rect 55180 40616 55338 40644
rect 55180 40604 55186 40616
rect 48961 40579 49019 40585
rect 48961 40545 48973 40579
rect 49007 40576 49019 40579
rect 49007 40548 49648 40576
rect 49007 40545 49019 40548
rect 48961 40539 49019 40545
rect 48041 40511 48099 40517
rect 44928 40480 47532 40508
rect 44928 40440 44956 40480
rect 41748 40412 42472 40440
rect 43640 40412 44956 40440
rect 41748 40400 41754 40412
rect 31726 40344 33180 40372
rect 33226 40332 33232 40384
rect 33284 40372 33290 40384
rect 34146 40372 34152 40384
rect 33284 40344 34152 40372
rect 33284 40332 33290 40344
rect 34146 40332 34152 40344
rect 34204 40332 34210 40384
rect 37090 40332 37096 40384
rect 37148 40372 37154 40384
rect 39942 40372 39948 40384
rect 37148 40344 39948 40372
rect 37148 40332 37154 40344
rect 39942 40332 39948 40344
rect 40000 40332 40006 40384
rect 40034 40332 40040 40384
rect 40092 40372 40098 40384
rect 40957 40375 41015 40381
rect 40957 40372 40969 40375
rect 40092 40344 40969 40372
rect 40092 40332 40098 40344
rect 40957 40341 40969 40344
rect 41003 40341 41015 40375
rect 40957 40335 41015 40341
rect 42058 40332 42064 40384
rect 42116 40372 42122 40384
rect 43640 40372 43668 40412
rect 47210 40400 47216 40452
rect 47268 40440 47274 40452
rect 47397 40443 47455 40449
rect 47397 40440 47409 40443
rect 47268 40412 47409 40440
rect 47268 40400 47274 40412
rect 47397 40409 47409 40412
rect 47443 40409 47455 40443
rect 47397 40403 47455 40409
rect 42116 40344 43668 40372
rect 42116 40332 42122 40344
rect 43714 40332 43720 40384
rect 43772 40372 43778 40384
rect 44085 40375 44143 40381
rect 44085 40372 44097 40375
rect 43772 40344 44097 40372
rect 43772 40332 43778 40344
rect 44085 40341 44097 40344
rect 44131 40341 44143 40375
rect 44085 40335 44143 40341
rect 45830 40332 45836 40384
rect 45888 40372 45894 40384
rect 46569 40375 46627 40381
rect 46569 40372 46581 40375
rect 45888 40344 46581 40372
rect 45888 40332 45894 40344
rect 46569 40341 46581 40344
rect 46615 40341 46627 40375
rect 47504 40372 47532 40480
rect 48041 40477 48053 40511
rect 48087 40477 48099 40511
rect 48041 40471 48099 40477
rect 49050 40468 49056 40520
rect 49108 40468 49114 40520
rect 49142 40468 49148 40520
rect 49200 40468 49206 40520
rect 49513 40511 49571 40517
rect 49513 40477 49525 40511
rect 49559 40477 49571 40511
rect 49513 40471 49571 40477
rect 47578 40400 47584 40452
rect 47636 40440 47642 40452
rect 49234 40440 49240 40452
rect 47636 40412 49240 40440
rect 47636 40400 47642 40412
rect 49234 40400 49240 40412
rect 49292 40440 49298 40452
rect 49528 40440 49556 40471
rect 49292 40412 49556 40440
rect 49292 40400 49298 40412
rect 48498 40372 48504 40384
rect 47504 40344 48504 40372
rect 46569 40335 46627 40341
rect 48498 40332 48504 40344
rect 48556 40332 48562 40384
rect 48590 40332 48596 40384
rect 48648 40332 48654 40384
rect 49620 40372 49648 40548
rect 49786 40536 49792 40588
rect 49844 40576 49850 40588
rect 50706 40576 50712 40588
rect 49844 40548 50712 40576
rect 49844 40536 49850 40548
rect 50706 40536 50712 40548
rect 50764 40536 50770 40588
rect 52178 40536 52184 40588
rect 52236 40536 52242 40588
rect 49697 40511 49755 40517
rect 49697 40477 49709 40511
rect 49743 40508 49755 40511
rect 50430 40508 50436 40520
rect 49743 40480 50436 40508
rect 49743 40477 49755 40480
rect 49697 40471 49755 40477
rect 50430 40468 50436 40480
rect 50488 40468 50494 40520
rect 53834 40468 53840 40520
rect 53892 40508 53898 40520
rect 53929 40511 53987 40517
rect 53929 40508 53941 40511
rect 53892 40480 53941 40508
rect 53892 40468 53898 40480
rect 53929 40477 53941 40480
rect 53975 40477 53987 40511
rect 53929 40471 53987 40477
rect 54570 40468 54576 40520
rect 54628 40468 54634 40520
rect 54849 40511 54907 40517
rect 54849 40477 54861 40511
rect 54895 40508 54907 40511
rect 55582 40508 55588 40520
rect 54895 40480 55588 40508
rect 54895 40477 54907 40480
rect 54849 40471 54907 40477
rect 55582 40468 55588 40480
rect 55640 40468 55646 40520
rect 56042 40468 56048 40520
rect 56100 40508 56106 40520
rect 56597 40511 56655 40517
rect 56597 40508 56609 40511
rect 56100 40480 56609 40508
rect 56100 40468 56106 40480
rect 56597 40477 56609 40480
rect 56643 40477 56655 40511
rect 56597 40471 56655 40477
rect 49878 40400 49884 40452
rect 49936 40440 49942 40452
rect 50157 40443 50215 40449
rect 50157 40440 50169 40443
rect 49936 40412 50169 40440
rect 49936 40400 49942 40412
rect 50157 40409 50169 40412
rect 50203 40409 50215 40443
rect 50157 40403 50215 40409
rect 51534 40400 51540 40452
rect 51592 40400 51598 40452
rect 50614 40372 50620 40384
rect 49620 40344 50620 40372
rect 50614 40332 50620 40344
rect 50672 40332 50678 40384
rect 52638 40332 52644 40384
rect 52696 40372 52702 40384
rect 53926 40372 53932 40384
rect 52696 40344 53932 40372
rect 52696 40332 52702 40344
rect 53926 40332 53932 40344
rect 53984 40372 53990 40384
rect 55030 40372 55036 40384
rect 53984 40344 55036 40372
rect 53984 40332 53990 40344
rect 55030 40332 55036 40344
rect 55088 40332 55094 40384
rect 552 40282 66424 40304
rect 552 40230 1998 40282
rect 2050 40230 2062 40282
rect 2114 40230 2126 40282
rect 2178 40230 2190 40282
rect 2242 40230 2254 40282
rect 2306 40230 49998 40282
rect 50050 40230 50062 40282
rect 50114 40230 50126 40282
rect 50178 40230 50190 40282
rect 50242 40230 50254 40282
rect 50306 40230 66424 40282
rect 552 40208 66424 40230
rect 8754 40128 8760 40180
rect 8812 40168 8818 40180
rect 10502 40168 10508 40180
rect 8812 40140 10508 40168
rect 8812 40128 8818 40140
rect 8570 40060 8576 40112
rect 8628 40100 8634 40112
rect 8628 40072 9352 40100
rect 8628 40060 8634 40072
rect 9324 40044 9352 40072
rect 9306 39992 9312 40044
rect 9364 39992 9370 40044
rect 9508 40041 9536 40140
rect 10502 40128 10508 40140
rect 10560 40128 10566 40180
rect 15215 40171 15273 40177
rect 15215 40137 15227 40171
rect 15261 40168 15273 40171
rect 15378 40168 15384 40180
rect 15261 40140 15384 40168
rect 15261 40137 15273 40140
rect 15215 40131 15273 40137
rect 15378 40128 15384 40140
rect 15436 40128 15442 40180
rect 17055 40171 17113 40177
rect 17055 40137 17067 40171
rect 17101 40168 17113 40171
rect 18690 40168 18696 40180
rect 17101 40140 18696 40168
rect 17101 40137 17113 40140
rect 17055 40131 17113 40137
rect 18690 40128 18696 40140
rect 18748 40128 18754 40180
rect 19324 40171 19382 40177
rect 19324 40137 19336 40171
rect 19370 40168 19382 40171
rect 19370 40140 20668 40168
rect 19370 40137 19382 40140
rect 19324 40131 19382 40137
rect 12526 40100 12532 40112
rect 12406 40072 12532 40100
rect 9493 40035 9551 40041
rect 9493 40001 9505 40035
rect 9539 40001 9551 40035
rect 9493 39995 9551 40001
rect 9769 40035 9827 40041
rect 9769 40001 9781 40035
rect 9815 40032 9827 40035
rect 10226 40032 10232 40044
rect 9815 40004 10232 40032
rect 9815 40001 9827 40004
rect 9769 39995 9827 40001
rect 10226 39992 10232 40004
rect 10284 39992 10290 40044
rect 10962 39992 10968 40044
rect 11020 39992 11026 40044
rect 11330 39992 11336 40044
rect 11388 40032 11394 40044
rect 11517 40035 11575 40041
rect 11517 40032 11529 40035
rect 11388 40004 11529 40032
rect 11388 39992 11394 40004
rect 11517 40001 11529 40004
rect 11563 40001 11575 40035
rect 11517 39995 11575 40001
rect 7650 39924 7656 39976
rect 7708 39924 7714 39976
rect 8205 39899 8263 39905
rect 8205 39865 8217 39899
rect 8251 39896 8263 39899
rect 9033 39899 9091 39905
rect 9033 39896 9045 39899
rect 8251 39868 9045 39896
rect 8251 39865 8263 39868
rect 8205 39859 8263 39865
rect 9033 39865 9045 39868
rect 9079 39865 9091 39899
rect 10980 39896 11008 39992
rect 12406 39896 12434 40072
rect 12526 40060 12532 40072
rect 12584 40060 12590 40112
rect 15470 40060 15476 40112
rect 15528 40060 15534 40112
rect 18322 40100 18328 40112
rect 18248 40072 18328 40100
rect 13722 39992 13728 40044
rect 13780 39992 13786 40044
rect 15488 40032 15516 40060
rect 15565 40035 15623 40041
rect 15565 40032 15577 40035
rect 15488 40004 15577 40032
rect 15565 40001 15577 40004
rect 15611 40032 15623 40035
rect 16482 40032 16488 40044
rect 15611 40004 16488 40032
rect 15611 40001 15623 40004
rect 15565 39995 15623 40001
rect 16482 39992 16488 40004
rect 16540 39992 16546 40044
rect 18248 40041 18276 40072
rect 18322 40060 18328 40072
rect 18380 40060 18386 40112
rect 20640 40100 20668 40140
rect 20714 40128 20720 40180
rect 20772 40168 20778 40180
rect 20901 40171 20959 40177
rect 20901 40168 20913 40171
rect 20772 40140 20913 40168
rect 20772 40128 20778 40140
rect 20901 40137 20913 40140
rect 20947 40137 20959 40171
rect 20901 40131 20959 40137
rect 21542 40128 21548 40180
rect 21600 40168 21606 40180
rect 21821 40171 21879 40177
rect 21821 40168 21833 40171
rect 21600 40140 21833 40168
rect 21600 40128 21606 40140
rect 21821 40137 21833 40140
rect 21867 40137 21879 40171
rect 21821 40131 21879 40137
rect 24844 40171 24902 40177
rect 24844 40137 24856 40171
rect 24890 40168 24902 40171
rect 25314 40168 25320 40180
rect 24890 40140 25320 40168
rect 24890 40137 24902 40140
rect 24844 40131 24902 40137
rect 25314 40128 25320 40140
rect 25372 40128 25378 40180
rect 27052 40171 27110 40177
rect 27052 40137 27064 40171
rect 27098 40168 27110 40171
rect 27430 40168 27436 40180
rect 27098 40140 27436 40168
rect 27098 40137 27110 40140
rect 27052 40131 27110 40137
rect 27430 40128 27436 40140
rect 27488 40128 27494 40180
rect 27522 40128 27528 40180
rect 27580 40168 27586 40180
rect 28537 40171 28595 40177
rect 27580 40140 28120 40168
rect 27580 40128 27586 40140
rect 21358 40100 21364 40112
rect 20640 40072 21364 40100
rect 21358 40060 21364 40072
rect 21416 40060 21422 40112
rect 21450 40060 21456 40112
rect 21508 40100 21514 40112
rect 22922 40100 22928 40112
rect 21508 40072 21588 40100
rect 21508 40060 21514 40072
rect 21560 40041 21588 40072
rect 22066 40072 22928 40100
rect 18233 40035 18291 40041
rect 18233 40001 18245 40035
rect 18279 40001 18291 40035
rect 21545 40035 21603 40041
rect 18233 39995 18291 40001
rect 20640 40004 21404 40032
rect 12805 39967 12863 39973
rect 12805 39933 12817 39967
rect 12851 39964 12863 39967
rect 12986 39964 12992 39976
rect 12851 39936 12992 39964
rect 12851 39933 12863 39936
rect 12805 39927 12863 39933
rect 12986 39924 12992 39936
rect 13044 39924 13050 39976
rect 15470 39924 15476 39976
rect 15528 39924 15534 39976
rect 17310 39924 17316 39976
rect 17368 39964 17374 39976
rect 19058 39964 19064 39976
rect 17368 39936 19064 39964
rect 17368 39924 17374 39936
rect 19058 39924 19064 39936
rect 19116 39924 19122 39976
rect 20438 39924 20444 39976
rect 20496 39924 20502 39976
rect 10980 39882 12434 39896
rect 10994 39868 12434 39882
rect 13357 39899 13415 39905
rect 9033 39859 9091 39865
rect 13357 39865 13369 39899
rect 13403 39896 13415 39899
rect 13906 39896 13912 39908
rect 13403 39868 13912 39896
rect 13403 39865 13415 39868
rect 13357 39859 13415 39865
rect 13906 39856 13912 39868
rect 13964 39856 13970 39908
rect 15746 39896 15752 39908
rect 14766 39868 15752 39896
rect 15746 39856 15752 39868
rect 15804 39896 15810 39908
rect 15804 39868 15870 39896
rect 16684 39868 18276 39896
rect 15804 39856 15810 39868
rect 8665 39831 8723 39837
rect 8665 39797 8677 39831
rect 8711 39828 8723 39831
rect 8846 39828 8852 39840
rect 8711 39800 8852 39828
rect 8711 39797 8723 39800
rect 8665 39791 8723 39797
rect 8846 39788 8852 39800
rect 8904 39788 8910 39840
rect 9122 39788 9128 39840
rect 9180 39788 9186 39840
rect 13078 39788 13084 39840
rect 13136 39828 13142 39840
rect 14182 39828 14188 39840
rect 13136 39800 14188 39828
rect 13136 39788 13142 39800
rect 14182 39788 14188 39800
rect 14240 39828 14246 39840
rect 16684 39828 16712 39868
rect 14240 39800 16712 39828
rect 14240 39788 14246 39800
rect 16942 39788 16948 39840
rect 17000 39828 17006 39840
rect 17589 39831 17647 39837
rect 17589 39828 17601 39831
rect 17000 39800 17601 39828
rect 17000 39788 17006 39800
rect 17589 39797 17601 39800
rect 17635 39797 17647 39831
rect 17589 39791 17647 39797
rect 17954 39788 17960 39840
rect 18012 39788 18018 39840
rect 18049 39831 18107 39837
rect 18049 39797 18061 39831
rect 18095 39828 18107 39831
rect 18138 39828 18144 39840
rect 18095 39800 18144 39828
rect 18095 39797 18107 39800
rect 18049 39791 18107 39797
rect 18138 39788 18144 39800
rect 18196 39788 18202 39840
rect 18248 39828 18276 39868
rect 20640 39828 20668 40004
rect 21266 39924 21272 39976
rect 21324 39924 21330 39976
rect 21376 39964 21404 40004
rect 21545 40001 21557 40035
rect 21591 40001 21603 40035
rect 21545 39995 21603 40001
rect 21818 39992 21824 40044
rect 21876 40032 21882 40044
rect 22066 40032 22094 40072
rect 21876 40004 22094 40032
rect 21876 39992 21882 40004
rect 22278 39992 22284 40044
rect 22336 39992 22342 40044
rect 22480 40041 22508 40072
rect 22922 40060 22928 40072
rect 22980 40060 22986 40112
rect 28092 40100 28120 40140
rect 28537 40137 28549 40171
rect 28583 40168 28595 40171
rect 29822 40168 29828 40180
rect 28583 40140 29828 40168
rect 28583 40137 28595 40140
rect 28537 40131 28595 40137
rect 29822 40128 29828 40140
rect 29880 40128 29886 40180
rect 29996 40171 30054 40177
rect 29996 40137 30008 40171
rect 30042 40168 30054 40171
rect 30650 40168 30656 40180
rect 30042 40140 30656 40168
rect 30042 40137 30054 40140
rect 29996 40131 30054 40137
rect 30650 40128 30656 40140
rect 30708 40128 30714 40180
rect 31478 40128 31484 40180
rect 31536 40128 31542 40180
rect 33042 40128 33048 40180
rect 33100 40177 33106 40180
rect 33100 40171 33115 40177
rect 33103 40137 33115 40171
rect 33100 40131 33115 40137
rect 33100 40128 33106 40131
rect 34054 40128 34060 40180
rect 34112 40168 34118 40180
rect 34149 40171 34207 40177
rect 34149 40168 34161 40171
rect 34112 40140 34161 40168
rect 34112 40128 34118 40140
rect 34149 40137 34161 40140
rect 34195 40137 34207 40171
rect 34149 40131 34207 40137
rect 35332 40171 35390 40177
rect 35332 40137 35344 40171
rect 35378 40168 35390 40171
rect 37458 40168 37464 40180
rect 35378 40140 37464 40168
rect 35378 40137 35390 40140
rect 35332 40131 35390 40137
rect 37458 40128 37464 40140
rect 37516 40128 37522 40180
rect 37632 40171 37690 40177
rect 37632 40137 37644 40171
rect 37678 40168 37690 40171
rect 38102 40168 38108 40180
rect 37678 40140 38108 40168
rect 37678 40137 37690 40140
rect 37632 40131 37690 40137
rect 38102 40128 38108 40140
rect 38160 40128 38166 40180
rect 39117 40171 39175 40177
rect 39117 40137 39129 40171
rect 39163 40168 39175 40171
rect 39666 40168 39672 40180
rect 39163 40140 39672 40168
rect 39163 40137 39175 40140
rect 39117 40131 39175 40137
rect 39666 40128 39672 40140
rect 39724 40128 39730 40180
rect 41414 40128 41420 40180
rect 41472 40168 41478 40180
rect 43257 40171 43315 40177
rect 41472 40140 42380 40168
rect 41472 40128 41478 40140
rect 28092 40072 28994 40100
rect 22465 40035 22523 40041
rect 22465 40001 22477 40035
rect 22511 40001 22523 40035
rect 22465 39995 22523 40001
rect 22646 39992 22652 40044
rect 22704 39992 22710 40044
rect 23290 39992 23296 40044
rect 23348 39992 23354 40044
rect 24581 40035 24639 40041
rect 24581 40001 24593 40035
rect 24627 40032 24639 40035
rect 26510 40032 26516 40044
rect 24627 40004 26516 40032
rect 24627 40001 24639 40004
rect 24581 39995 24639 40001
rect 26510 39992 26516 40004
rect 26568 40032 26574 40044
rect 27154 40032 27160 40044
rect 26568 40004 27160 40032
rect 26568 39992 26574 40004
rect 27154 39992 27160 40004
rect 27212 39992 27218 40044
rect 28966 40032 28994 40072
rect 33502 40060 33508 40112
rect 33560 40100 33566 40112
rect 34514 40100 34520 40112
rect 33560 40072 34520 40100
rect 33560 40060 33566 40072
rect 34514 40060 34520 40072
rect 34572 40060 34578 40112
rect 34974 40100 34980 40112
rect 34716 40072 34980 40100
rect 31846 40032 31852 40044
rect 28966 40004 31852 40032
rect 31846 39992 31852 40004
rect 31904 39992 31910 40044
rect 32582 40032 32588 40044
rect 32048 40004 32588 40032
rect 23474 39964 23480 39976
rect 21376 39936 23480 39964
rect 23474 39924 23480 39936
rect 23532 39924 23538 39976
rect 24026 39924 24032 39976
rect 24084 39964 24090 39976
rect 24397 39967 24455 39973
rect 24397 39964 24409 39967
rect 24084 39936 24409 39964
rect 24084 39924 24090 39936
rect 24397 39933 24409 39936
rect 24443 39933 24455 39967
rect 24397 39927 24455 39933
rect 26234 39924 26240 39976
rect 26292 39964 26298 39976
rect 26789 39967 26847 39973
rect 26789 39964 26801 39967
rect 26292 39936 26801 39964
rect 26292 39924 26298 39936
rect 26789 39933 26801 39936
rect 26835 39933 26847 39967
rect 26789 39927 26847 39933
rect 29546 39924 29552 39976
rect 29604 39964 29610 39976
rect 29733 39967 29791 39973
rect 29733 39964 29745 39967
rect 29604 39936 29745 39964
rect 29604 39924 29610 39936
rect 29733 39933 29745 39936
rect 29779 39933 29791 39967
rect 32048 39964 32076 40004
rect 32582 39992 32588 40004
rect 32640 39992 32646 40044
rect 34716 40041 34744 40072
rect 34974 40060 34980 40072
rect 35032 40060 35038 40112
rect 39390 40060 39396 40112
rect 39448 40100 39454 40112
rect 39448 40072 39804 40100
rect 39448 40060 39454 40072
rect 34701 40035 34759 40041
rect 34701 40001 34713 40035
rect 34747 40001 34759 40035
rect 34701 39995 34759 40001
rect 36817 40035 36875 40041
rect 36817 40001 36829 40035
rect 36863 40032 36875 40035
rect 37274 40032 37280 40044
rect 36863 40004 37280 40032
rect 36863 40001 36875 40004
rect 36817 39995 36875 40001
rect 37274 39992 37280 40004
rect 37332 39992 37338 40044
rect 37366 39992 37372 40044
rect 37424 39992 37430 40044
rect 38654 39992 38660 40044
rect 38712 40032 38718 40044
rect 39776 40032 39804 40072
rect 41598 40060 41604 40112
rect 41656 40100 41662 40112
rect 42352 40100 42380 40140
rect 43257 40137 43269 40171
rect 43303 40168 43315 40171
rect 43346 40168 43352 40180
rect 43303 40140 43352 40168
rect 43303 40137 43315 40140
rect 43257 40131 43315 40137
rect 43346 40128 43352 40140
rect 43404 40128 43410 40180
rect 45738 40128 45744 40180
rect 45796 40168 45802 40180
rect 46569 40171 46627 40177
rect 46569 40168 46581 40171
rect 45796 40140 46581 40168
rect 45796 40128 45802 40140
rect 46569 40137 46581 40140
rect 46615 40137 46627 40171
rect 46569 40131 46627 40137
rect 47936 40171 47994 40177
rect 47936 40137 47948 40171
rect 47982 40168 47994 40171
rect 48590 40168 48596 40180
rect 47982 40140 48596 40168
rect 47982 40137 47994 40140
rect 47936 40131 47994 40137
rect 43806 40100 43812 40112
rect 41656 40072 42012 40100
rect 41656 40060 41662 40072
rect 38712 40004 39712 40032
rect 39776 40004 41460 40032
rect 38712 39992 38718 40004
rect 31142 39936 32076 39964
rect 33321 39967 33379 39973
rect 29733 39927 29791 39933
rect 33321 39933 33333 39967
rect 33367 39964 33379 39967
rect 33367 39936 34836 39964
rect 33367 39933 33379 39936
rect 33321 39927 33379 39933
rect 21726 39896 21732 39908
rect 20824 39868 21732 39896
rect 20824 39837 20852 39868
rect 21726 39856 21732 39868
rect 21784 39856 21790 39908
rect 22189 39899 22247 39905
rect 22189 39865 22201 39899
rect 22235 39896 22247 39899
rect 24854 39896 24860 39908
rect 22235 39868 24860 39896
rect 22235 39865 22247 39868
rect 22189 39859 22247 39865
rect 24854 39856 24860 39868
rect 24912 39856 24918 39908
rect 24946 39856 24952 39908
rect 25004 39896 25010 39908
rect 25004 39868 25346 39896
rect 26160 39868 27554 39896
rect 25004 39856 25010 39868
rect 18248 39800 20668 39828
rect 20809 39831 20867 39837
rect 20809 39797 20821 39831
rect 20855 39797 20867 39831
rect 20809 39791 20867 39797
rect 21266 39788 21272 39840
rect 21324 39828 21330 39840
rect 21361 39831 21419 39837
rect 21361 39828 21373 39831
rect 21324 39800 21373 39828
rect 21324 39788 21330 39800
rect 21361 39797 21373 39800
rect 21407 39797 21419 39831
rect 21361 39791 21419 39797
rect 23842 39788 23848 39840
rect 23900 39788 23906 39840
rect 25240 39828 25268 39868
rect 26160 39828 26188 39868
rect 32582 39856 32588 39908
rect 32640 39896 32646 39908
rect 32950 39896 32956 39908
rect 32640 39868 32956 39896
rect 32640 39856 32646 39868
rect 32950 39856 32956 39868
rect 33008 39856 33014 39908
rect 33778 39856 33784 39908
rect 33836 39896 33842 39908
rect 34517 39899 34575 39905
rect 34517 39896 34529 39899
rect 33836 39868 34529 39896
rect 33836 39856 33842 39868
rect 34517 39865 34529 39868
rect 34563 39865 34575 39899
rect 34808 39896 34836 39936
rect 34882 39924 34888 39976
rect 34940 39964 34946 39976
rect 35069 39967 35127 39973
rect 35069 39964 35081 39967
rect 34940 39936 35081 39964
rect 34940 39924 34946 39936
rect 35069 39933 35081 39936
rect 35115 39933 35127 39967
rect 39684 39964 39712 40004
rect 39758 39964 39764 39976
rect 39684 39936 39764 39964
rect 35069 39927 35127 39933
rect 39758 39924 39764 39936
rect 39816 39924 39822 39976
rect 41046 39924 41052 39976
rect 41104 39964 41110 39976
rect 41104 39936 41170 39964
rect 41104 39924 41110 39936
rect 35618 39896 35624 39908
rect 34808 39868 35624 39896
rect 34517 39859 34575 39865
rect 35618 39856 35624 39868
rect 35676 39856 35682 39908
rect 36078 39856 36084 39908
rect 36136 39856 36142 39908
rect 38102 39856 38108 39908
rect 38160 39856 38166 39908
rect 40034 39856 40040 39908
rect 40092 39856 40098 39908
rect 41432 39896 41460 40004
rect 41984 39973 42012 40072
rect 42352 40072 43812 40100
rect 42245 40035 42303 40041
rect 42245 40001 42257 40035
rect 42291 40032 42303 40035
rect 42352 40032 42380 40072
rect 43806 40060 43812 40072
rect 43864 40060 43870 40112
rect 43990 40100 43996 40112
rect 43916 40072 43996 40100
rect 42291 40004 42380 40032
rect 42291 40001 42303 40004
rect 42245 39995 42303 40001
rect 43070 39992 43076 40044
rect 43128 40032 43134 40044
rect 43530 40032 43536 40044
rect 43128 40004 43536 40032
rect 43128 39992 43134 40004
rect 43530 39992 43536 40004
rect 43588 39992 43594 40044
rect 43916 40041 43944 40072
rect 43990 40060 43996 40072
rect 44048 40060 44054 40112
rect 43901 40035 43959 40041
rect 43901 40001 43913 40035
rect 43947 40001 43959 40035
rect 43901 39995 43959 40001
rect 44818 39992 44824 40044
rect 44876 39992 44882 40044
rect 45097 40035 45155 40041
rect 45097 40001 45109 40035
rect 45143 40032 45155 40035
rect 46106 40032 46112 40044
rect 45143 40004 46112 40032
rect 45143 40001 45155 40004
rect 45097 39995 45155 40001
rect 46106 39992 46112 40004
rect 46164 39992 46170 40044
rect 46584 40032 46612 40131
rect 48590 40128 48596 40140
rect 48648 40128 48654 40180
rect 49602 40168 49608 40180
rect 49252 40140 49608 40168
rect 47213 40035 47271 40041
rect 47213 40032 47225 40035
rect 46584 40004 47225 40032
rect 47213 40001 47225 40004
rect 47259 40001 47271 40035
rect 47213 39995 47271 40001
rect 47673 40035 47731 40041
rect 47673 40001 47685 40035
rect 47719 40032 47731 40035
rect 49252 40032 49280 40140
rect 49602 40128 49608 40140
rect 49660 40168 49666 40180
rect 51350 40168 51356 40180
rect 49660 40140 51356 40168
rect 49660 40128 49666 40140
rect 51350 40128 51356 40140
rect 51408 40128 51414 40180
rect 54570 40168 54576 40180
rect 51552 40140 54576 40168
rect 51552 40112 51580 40140
rect 49878 40060 49884 40112
rect 49936 40100 49942 40112
rect 50430 40100 50436 40112
rect 49936 40072 50436 40100
rect 49936 40060 49942 40072
rect 50430 40060 50436 40072
rect 50488 40060 50494 40112
rect 51534 40100 51540 40112
rect 51046 40072 51540 40100
rect 47719 40004 49280 40032
rect 47719 40001 47731 40004
rect 47673 39995 47731 40001
rect 49694 39992 49700 40044
rect 49752 39992 49758 40044
rect 41969 39967 42027 39973
rect 41969 39933 41981 39967
rect 42015 39964 42027 39967
rect 42150 39964 42156 39976
rect 42015 39936 42156 39964
rect 42015 39933 42027 39936
rect 41969 39927 42027 39933
rect 42150 39924 42156 39936
rect 42208 39924 42214 39976
rect 49712 39936 50660 39964
rect 46474 39896 46480 39908
rect 41432 39868 43852 39896
rect 46322 39868 46480 39896
rect 25240 39800 26188 39828
rect 26326 39788 26332 39840
rect 26384 39828 26390 39840
rect 27062 39828 27068 39840
rect 26384 39800 27068 39828
rect 26384 39788 26390 39800
rect 27062 39788 27068 39800
rect 27120 39828 27126 39840
rect 27430 39828 27436 39840
rect 27120 39800 27436 39828
rect 27120 39788 27126 39800
rect 27430 39788 27436 39800
rect 27488 39788 27494 39840
rect 28350 39788 28356 39840
rect 28408 39828 28414 39840
rect 31018 39828 31024 39840
rect 28408 39800 31024 39828
rect 28408 39788 28414 39800
rect 31018 39788 31024 39800
rect 31076 39788 31082 39840
rect 31573 39831 31631 39837
rect 31573 39797 31585 39831
rect 31619 39828 31631 39831
rect 33796 39828 33824 39856
rect 31619 39800 33824 39828
rect 34609 39831 34667 39837
rect 31619 39797 31631 39800
rect 31573 39791 31631 39797
rect 34609 39797 34621 39831
rect 34655 39828 34667 39831
rect 41046 39828 41052 39840
rect 34655 39800 41052 39828
rect 34655 39797 34667 39800
rect 34609 39791 34667 39797
rect 41046 39788 41052 39800
rect 41104 39788 41110 39840
rect 41506 39788 41512 39840
rect 41564 39788 41570 39840
rect 41598 39788 41604 39840
rect 41656 39788 41662 39840
rect 41966 39788 41972 39840
rect 42024 39828 42030 39840
rect 42061 39831 42119 39837
rect 42061 39828 42073 39831
rect 42024 39800 42073 39828
rect 42024 39788 42030 39800
rect 42061 39797 42073 39800
rect 42107 39797 42119 39831
rect 42061 39791 42119 39797
rect 43530 39788 43536 39840
rect 43588 39828 43594 39840
rect 43625 39831 43683 39837
rect 43625 39828 43637 39831
rect 43588 39800 43637 39828
rect 43588 39788 43594 39800
rect 43625 39797 43637 39800
rect 43671 39797 43683 39831
rect 43625 39791 43683 39797
rect 43714 39788 43720 39840
rect 43772 39788 43778 39840
rect 43824 39828 43852 39868
rect 46474 39856 46480 39868
rect 46532 39856 46538 39908
rect 46584 39868 48314 39896
rect 46584 39828 46612 39868
rect 43824 39800 46612 39828
rect 46658 39788 46664 39840
rect 46716 39788 46722 39840
rect 48286 39828 48314 39868
rect 48958 39856 48964 39908
rect 49016 39856 49022 39908
rect 49712 39896 49740 39936
rect 49252 39868 49740 39896
rect 49804 39868 50016 39896
rect 49252 39828 49280 39868
rect 48286 39800 49280 39828
rect 49421 39831 49479 39837
rect 49421 39797 49433 39831
rect 49467 39828 49479 39831
rect 49804 39828 49832 39868
rect 49988 39840 50016 39868
rect 49467 39800 49832 39828
rect 49467 39797 49479 39800
rect 49421 39791 49479 39797
rect 49878 39788 49884 39840
rect 49936 39788 49942 39840
rect 49970 39788 49976 39840
rect 50028 39788 50034 39840
rect 50246 39788 50252 39840
rect 50304 39828 50310 39840
rect 50341 39831 50399 39837
rect 50341 39828 50353 39831
rect 50304 39800 50353 39828
rect 50304 39788 50310 39800
rect 50341 39797 50353 39800
rect 50387 39797 50399 39831
rect 50632 39828 50660 39936
rect 50706 39856 50712 39908
rect 50764 39896 50770 39908
rect 51046 39896 51074 40072
rect 51534 40060 51540 40072
rect 51592 40060 51598 40112
rect 53466 39992 53472 40044
rect 53524 40032 53530 40044
rect 54128 40041 54156 40140
rect 54570 40128 54576 40140
rect 54628 40128 54634 40180
rect 55582 40128 55588 40180
rect 55640 40128 55646 40180
rect 55030 40060 55036 40112
rect 55088 40060 55094 40112
rect 60734 40060 60740 40112
rect 60792 40100 60798 40112
rect 64966 40100 64972 40112
rect 60792 40072 64972 40100
rect 60792 40060 60798 40072
rect 64966 40060 64972 40072
rect 65024 40060 65030 40112
rect 53837 40035 53895 40041
rect 53837 40032 53849 40035
rect 53524 40004 53849 40032
rect 53524 39992 53530 40004
rect 53837 40001 53849 40004
rect 53883 40001 53895 40035
rect 53837 39995 53895 40001
rect 54113 40035 54171 40041
rect 54113 40001 54125 40035
rect 54159 40001 54171 40035
rect 54113 39995 54171 40001
rect 54662 39992 54668 40044
rect 54720 40032 54726 40044
rect 54849 40035 54907 40041
rect 54849 40032 54861 40035
rect 54720 40004 54861 40032
rect 54720 39992 54726 40004
rect 54849 40001 54861 40004
rect 54895 40001 54907 40035
rect 54849 39995 54907 40001
rect 55048 39973 55076 40060
rect 56226 39992 56232 40044
rect 56284 39992 56290 40044
rect 55033 39967 55091 39973
rect 55033 39933 55045 39967
rect 55079 39933 55091 39967
rect 55033 39927 55091 39933
rect 55953 39967 56011 39973
rect 55953 39933 55965 39967
rect 55999 39964 56011 39967
rect 56502 39964 56508 39976
rect 55999 39936 56508 39964
rect 55999 39933 56011 39936
rect 55953 39927 56011 39933
rect 56502 39924 56508 39936
rect 56560 39924 56566 39976
rect 50764 39868 51074 39896
rect 50764 39856 50770 39868
rect 52086 39856 52092 39908
rect 52144 39856 52150 39908
rect 53098 39856 53104 39908
rect 53156 39856 53162 39908
rect 56042 39896 56048 39908
rect 55140 39868 56048 39896
rect 52822 39828 52828 39840
rect 50632 39800 52828 39828
rect 50341 39791 50399 39797
rect 52822 39788 52828 39800
rect 52880 39788 52886 39840
rect 54478 39788 54484 39840
rect 54536 39828 54542 39840
rect 55140 39837 55168 39868
rect 56042 39856 56048 39868
rect 56100 39856 56106 39908
rect 55125 39831 55183 39837
rect 55125 39828 55137 39831
rect 54536 39800 55137 39828
rect 54536 39788 54542 39800
rect 55125 39797 55137 39800
rect 55171 39797 55183 39831
rect 55125 39791 55183 39797
rect 55306 39788 55312 39840
rect 55364 39828 55370 39840
rect 55493 39831 55551 39837
rect 55493 39828 55505 39831
rect 55364 39800 55505 39828
rect 55364 39788 55370 39800
rect 55493 39797 55505 39800
rect 55539 39797 55551 39831
rect 55493 39791 55551 39797
rect 552 39738 66424 39760
rect 552 39686 2918 39738
rect 2970 39686 2982 39738
rect 3034 39686 3046 39738
rect 3098 39686 3110 39738
rect 3162 39686 3174 39738
rect 3226 39686 50918 39738
rect 50970 39686 50982 39738
rect 51034 39686 51046 39738
rect 51098 39686 51110 39738
rect 51162 39686 51174 39738
rect 51226 39686 66424 39738
rect 552 39664 66424 39686
rect 12802 39624 12808 39636
rect 9140 39596 12808 39624
rect 8570 39556 8576 39568
rect 8418 39528 8576 39556
rect 8570 39516 8576 39528
rect 8628 39516 8634 39568
rect 8846 39516 8852 39568
rect 8904 39516 8910 39568
rect 9140 39497 9168 39596
rect 12802 39584 12808 39596
rect 12860 39624 12866 39636
rect 17310 39624 17316 39636
rect 12860 39596 17316 39624
rect 12860 39584 12866 39596
rect 9490 39516 9496 39568
rect 9548 39556 9554 39568
rect 9677 39559 9735 39565
rect 9677 39556 9689 39559
rect 9548 39528 9689 39556
rect 9548 39516 9554 39528
rect 9677 39525 9689 39528
rect 9723 39556 9735 39559
rect 11422 39556 11428 39568
rect 9723 39528 11428 39556
rect 9723 39525 9735 39528
rect 9677 39519 9735 39525
rect 11422 39516 11428 39528
rect 11480 39516 11486 39568
rect 12434 39516 12440 39568
rect 12492 39516 12498 39568
rect 13538 39516 13544 39568
rect 13596 39556 13602 39568
rect 15470 39556 15476 39568
rect 13596 39528 15476 39556
rect 13596 39516 13602 39528
rect 9125 39491 9183 39497
rect 9125 39457 9137 39491
rect 9171 39457 9183 39491
rect 9125 39451 9183 39457
rect 9585 39491 9643 39497
rect 9585 39457 9597 39491
rect 9631 39457 9643 39491
rect 9585 39451 9643 39457
rect 11333 39491 11391 39497
rect 11333 39457 11345 39491
rect 11379 39488 11391 39491
rect 11698 39488 11704 39500
rect 11379 39460 11704 39488
rect 11379 39457 11391 39460
rect 11333 39451 11391 39457
rect 7377 39423 7435 39429
rect 7377 39389 7389 39423
rect 7423 39420 7435 39423
rect 7650 39420 7656 39432
rect 7423 39392 7656 39420
rect 7423 39389 7435 39392
rect 7377 39383 7435 39389
rect 7650 39380 7656 39392
rect 7708 39420 7714 39432
rect 9600 39420 9628 39451
rect 11698 39448 11704 39460
rect 11756 39448 11762 39500
rect 13740 39497 13768 39528
rect 15470 39516 15476 39528
rect 15528 39516 15534 39568
rect 15562 39516 15568 39568
rect 15620 39516 15626 39568
rect 13725 39491 13783 39497
rect 13725 39457 13737 39491
rect 13771 39457 13783 39491
rect 13725 39451 13783 39457
rect 13906 39448 13912 39500
rect 13964 39488 13970 39500
rect 14185 39491 14243 39497
rect 14185 39488 14197 39491
rect 13964 39460 14197 39488
rect 13964 39448 13970 39460
rect 14185 39457 14197 39460
rect 14231 39457 14243 39491
rect 14185 39451 14243 39457
rect 14277 39491 14335 39497
rect 14277 39457 14289 39491
rect 14323 39488 14335 39491
rect 14458 39488 14464 39500
rect 14323 39460 14464 39488
rect 14323 39457 14335 39460
rect 14277 39451 14335 39457
rect 14458 39448 14464 39460
rect 14516 39448 14522 39500
rect 16684 39497 16712 39596
rect 17310 39584 17316 39596
rect 17368 39584 17374 39636
rect 18414 39584 18420 39636
rect 18472 39584 18478 39636
rect 19058 39584 19064 39636
rect 19116 39624 19122 39636
rect 20441 39627 20499 39633
rect 20441 39624 20453 39627
rect 19116 39596 20453 39624
rect 19116 39584 19122 39596
rect 20441 39593 20453 39596
rect 20487 39593 20499 39627
rect 20441 39587 20499 39593
rect 21266 39584 21272 39636
rect 21324 39584 21330 39636
rect 21358 39584 21364 39636
rect 21416 39624 21422 39636
rect 22097 39627 22155 39633
rect 22097 39624 22109 39627
rect 21416 39596 22109 39624
rect 21416 39584 21422 39596
rect 22097 39593 22109 39596
rect 22143 39593 22155 39627
rect 22097 39587 22155 39593
rect 22465 39627 22523 39633
rect 22465 39593 22477 39627
rect 22511 39624 22523 39627
rect 22738 39624 22744 39636
rect 22511 39596 22744 39624
rect 22511 39593 22523 39596
rect 22465 39587 22523 39593
rect 22738 39584 22744 39596
rect 22796 39584 22802 39636
rect 24026 39584 24032 39636
rect 24084 39584 24090 39636
rect 25130 39584 25136 39636
rect 25188 39584 25194 39636
rect 25501 39627 25559 39633
rect 25501 39593 25513 39627
rect 25547 39624 25559 39627
rect 26326 39624 26332 39636
rect 25547 39596 26332 39624
rect 25547 39593 25559 39596
rect 25501 39587 25559 39593
rect 26326 39584 26332 39596
rect 26384 39584 26390 39636
rect 28350 39624 28356 39636
rect 27540 39596 28356 39624
rect 16942 39516 16948 39568
rect 17000 39516 17006 39568
rect 18506 39516 18512 39568
rect 18564 39556 18570 39568
rect 19153 39559 19211 39565
rect 19153 39556 19165 39559
rect 18564 39528 19165 39556
rect 18564 39516 18570 39528
rect 19153 39525 19165 39528
rect 19199 39556 19211 39559
rect 24670 39556 24676 39568
rect 19199 39528 24676 39556
rect 19199 39525 19211 39528
rect 19153 39519 19211 39525
rect 24670 39516 24676 39528
rect 24728 39516 24734 39568
rect 24854 39516 24860 39568
rect 24912 39556 24918 39568
rect 27540 39556 27568 39596
rect 28350 39584 28356 39596
rect 28408 39584 28414 39636
rect 28445 39627 28503 39633
rect 28445 39593 28457 39627
rect 28491 39624 28503 39627
rect 28718 39624 28724 39636
rect 28491 39596 28724 39624
rect 28491 39593 28503 39596
rect 28445 39587 28503 39593
rect 28718 39584 28724 39596
rect 28776 39584 28782 39636
rect 28813 39627 28871 39633
rect 28813 39593 28825 39627
rect 28859 39624 28871 39627
rect 29362 39624 29368 39636
rect 28859 39596 29368 39624
rect 28859 39593 28871 39596
rect 28813 39587 28871 39593
rect 29362 39584 29368 39596
rect 29420 39584 29426 39636
rect 31021 39627 31079 39633
rect 31021 39593 31033 39627
rect 31067 39624 31079 39627
rect 31478 39624 31484 39636
rect 31067 39596 31484 39624
rect 31067 39593 31079 39596
rect 31021 39587 31079 39593
rect 31478 39584 31484 39596
rect 31536 39584 31542 39636
rect 33226 39624 33232 39636
rect 32232 39596 33232 39624
rect 24912 39528 27568 39556
rect 24912 39516 24918 39528
rect 27614 39516 27620 39568
rect 27672 39556 27678 39568
rect 30374 39556 30380 39568
rect 27672 39528 30380 39556
rect 27672 39516 27678 39528
rect 30374 39516 30380 39528
rect 30432 39516 30438 39568
rect 32232 39556 32260 39596
rect 33226 39584 33232 39596
rect 33284 39584 33290 39636
rect 33413 39627 33471 39633
rect 33413 39593 33425 39627
rect 33459 39624 33471 39627
rect 33594 39624 33600 39636
rect 33459 39596 33600 39624
rect 33459 39593 33471 39596
rect 33413 39587 33471 39593
rect 33594 39584 33600 39596
rect 33652 39584 33658 39636
rect 33686 39584 33692 39636
rect 33744 39624 33750 39636
rect 33873 39627 33931 39633
rect 33873 39624 33885 39627
rect 33744 39596 33885 39624
rect 33744 39584 33750 39596
rect 33873 39593 33885 39596
rect 33919 39593 33931 39627
rect 33873 39587 33931 39593
rect 34606 39584 34612 39636
rect 34664 39624 34670 39636
rect 35250 39624 35256 39636
rect 34664 39596 35256 39624
rect 34664 39584 34670 39596
rect 35250 39584 35256 39596
rect 35308 39584 35314 39636
rect 35986 39584 35992 39636
rect 36044 39624 36050 39636
rect 36081 39627 36139 39633
rect 36081 39624 36093 39627
rect 36044 39596 36093 39624
rect 36044 39584 36050 39596
rect 36081 39593 36093 39596
rect 36127 39593 36139 39627
rect 36081 39587 36139 39593
rect 36541 39627 36599 39633
rect 36541 39593 36553 39627
rect 36587 39624 36599 39627
rect 36587 39596 38332 39624
rect 36587 39593 36599 39596
rect 36541 39587 36599 39593
rect 31496 39528 32260 39556
rect 16669 39491 16727 39497
rect 16669 39457 16681 39491
rect 16715 39457 16727 39491
rect 16669 39451 16727 39457
rect 18046 39448 18052 39500
rect 18104 39448 18110 39500
rect 21542 39448 21548 39500
rect 21600 39488 21606 39500
rect 21637 39491 21695 39497
rect 21637 39488 21649 39491
rect 21600 39460 21649 39488
rect 21600 39448 21606 39460
rect 21637 39457 21649 39460
rect 21683 39457 21695 39491
rect 21637 39451 21695 39457
rect 21726 39448 21732 39500
rect 21784 39448 21790 39500
rect 28718 39488 28724 39500
rect 25792 39460 28724 39488
rect 7708 39392 9628 39420
rect 9769 39423 9827 39429
rect 7708 39380 7714 39392
rect 9769 39389 9781 39423
rect 9815 39389 9827 39423
rect 9769 39383 9827 39389
rect 11609 39423 11667 39429
rect 11609 39389 11621 39423
rect 11655 39420 11667 39423
rect 13078 39420 13084 39432
rect 11655 39392 13084 39420
rect 11655 39389 11667 39392
rect 11609 39383 11667 39389
rect 9582 39312 9588 39364
rect 9640 39352 9646 39364
rect 9784 39352 9812 39383
rect 13078 39380 13084 39392
rect 13136 39380 13142 39432
rect 13449 39423 13507 39429
rect 13449 39389 13461 39423
rect 13495 39420 13507 39423
rect 13495 39392 13860 39420
rect 13495 39389 13507 39392
rect 13449 39383 13507 39389
rect 9640 39324 9812 39352
rect 9640 39312 9646 39324
rect 10410 39312 10416 39364
rect 10468 39352 10474 39364
rect 13832 39361 13860 39392
rect 14366 39380 14372 39432
rect 14424 39380 14430 39432
rect 15286 39380 15292 39432
rect 15344 39380 15350 39432
rect 15473 39423 15531 39429
rect 15473 39389 15485 39423
rect 15519 39420 15531 39423
rect 17402 39420 17408 39432
rect 15519 39392 17408 39420
rect 15519 39389 15531 39392
rect 15473 39383 15531 39389
rect 17402 39380 17408 39392
rect 17460 39380 17466 39432
rect 20806 39380 20812 39432
rect 20864 39420 20870 39432
rect 21818 39420 21824 39432
rect 20864 39392 21824 39420
rect 20864 39380 20870 39392
rect 21818 39380 21824 39392
rect 21876 39380 21882 39432
rect 22557 39423 22615 39429
rect 22557 39420 22569 39423
rect 22066 39392 22569 39420
rect 10965 39355 11023 39361
rect 10965 39352 10977 39355
rect 10468 39324 10977 39352
rect 10468 39312 10474 39324
rect 10965 39321 10977 39324
rect 11011 39321 11023 39355
rect 10965 39315 11023 39321
rect 13817 39355 13875 39361
rect 13817 39321 13829 39355
rect 13863 39321 13875 39355
rect 13817 39315 13875 39321
rect 15930 39312 15936 39364
rect 15988 39312 15994 39364
rect 8846 39244 8852 39296
rect 8904 39284 8910 39296
rect 9217 39287 9275 39293
rect 9217 39284 9229 39287
rect 8904 39256 9229 39284
rect 8904 39244 8910 39256
rect 9217 39253 9229 39256
rect 9263 39253 9275 39287
rect 9217 39247 9275 39253
rect 11977 39287 12035 39293
rect 11977 39253 11989 39287
rect 12023 39284 12035 39287
rect 12986 39284 12992 39296
rect 12023 39256 12992 39284
rect 12023 39253 12035 39256
rect 11977 39247 12035 39253
rect 12986 39244 12992 39256
rect 13044 39244 13050 39296
rect 20530 39244 20536 39296
rect 20588 39284 20594 39296
rect 22066 39284 22094 39392
rect 22557 39389 22569 39392
rect 22603 39389 22615 39423
rect 22557 39383 22615 39389
rect 22646 39380 22652 39432
rect 22704 39380 22710 39432
rect 23845 39423 23903 39429
rect 23845 39389 23857 39423
rect 23891 39389 23903 39423
rect 23845 39383 23903 39389
rect 23937 39423 23995 39429
rect 23937 39389 23949 39423
rect 23983 39420 23995 39423
rect 24302 39420 24308 39432
rect 23983 39392 24308 39420
rect 23983 39389 23995 39392
rect 23937 39383 23995 39389
rect 22462 39312 22468 39364
rect 22520 39352 22526 39364
rect 23860 39352 23888 39383
rect 24302 39380 24308 39392
rect 24360 39380 24366 39432
rect 25590 39380 25596 39432
rect 25648 39380 25654 39432
rect 25792 39429 25820 39460
rect 28718 39448 28724 39460
rect 28776 39448 28782 39500
rect 29825 39491 29883 39497
rect 29825 39488 29837 39491
rect 28920 39460 29837 39488
rect 25777 39423 25835 39429
rect 25777 39389 25789 39423
rect 25823 39389 25835 39423
rect 25777 39383 25835 39389
rect 26418 39380 26424 39432
rect 26476 39420 26482 39432
rect 26973 39423 27031 39429
rect 26973 39420 26985 39423
rect 26476 39392 26985 39420
rect 26476 39380 26482 39392
rect 26973 39389 26985 39392
rect 27019 39389 27031 39423
rect 26973 39383 27031 39389
rect 27709 39423 27767 39429
rect 27709 39389 27721 39423
rect 27755 39389 27767 39423
rect 27709 39383 27767 39389
rect 26050 39352 26056 39364
rect 22520 39324 26056 39352
rect 22520 39312 22526 39324
rect 26050 39312 26056 39324
rect 26108 39312 26114 39364
rect 27614 39312 27620 39364
rect 27672 39352 27678 39364
rect 27724 39352 27752 39383
rect 28810 39380 28816 39432
rect 28868 39420 28874 39432
rect 28920 39429 28948 39460
rect 29825 39457 29837 39460
rect 29871 39457 29883 39491
rect 31496 39488 31524 39528
rect 34514 39516 34520 39568
rect 34572 39556 34578 39568
rect 36173 39559 36231 39565
rect 34572 39528 35940 39556
rect 34572 39516 34578 39528
rect 29825 39451 29883 39457
rect 30024 39460 31524 39488
rect 28905 39423 28963 39429
rect 28905 39420 28917 39423
rect 28868 39392 28917 39420
rect 28868 39380 28874 39392
rect 28905 39389 28917 39392
rect 28951 39389 28963 39423
rect 28905 39383 28963 39389
rect 28994 39380 29000 39432
rect 29052 39380 29058 39432
rect 27672 39324 27752 39352
rect 27672 39312 27678 39324
rect 27890 39312 27896 39364
rect 27948 39352 27954 39364
rect 30024 39352 30052 39460
rect 31570 39448 31576 39500
rect 31628 39448 31634 39500
rect 32950 39448 32956 39500
rect 33008 39448 33014 39500
rect 33410 39448 33416 39500
rect 33468 39488 33474 39500
rect 33781 39491 33839 39497
rect 33781 39488 33793 39491
rect 33468 39460 33793 39488
rect 33468 39448 33474 39460
rect 33781 39457 33793 39460
rect 33827 39457 33839 39491
rect 35912 39488 35940 39528
rect 36173 39525 36185 39559
rect 36219 39556 36231 39559
rect 36630 39556 36636 39568
rect 36219 39528 36636 39556
rect 36219 39525 36231 39528
rect 36173 39519 36231 39525
rect 36630 39516 36636 39528
rect 36688 39516 36694 39568
rect 36998 39516 37004 39568
rect 37056 39516 37062 39568
rect 38304 39556 38332 39596
rect 38562 39584 38568 39636
rect 38620 39584 38626 39636
rect 38930 39584 38936 39636
rect 38988 39584 38994 39636
rect 42889 39627 42947 39633
rect 42889 39624 42901 39627
rect 40052 39596 41092 39624
rect 39025 39559 39083 39565
rect 39025 39556 39037 39559
rect 38304 39528 39037 39556
rect 39025 39525 39037 39528
rect 39071 39525 39083 39559
rect 39025 39519 39083 39525
rect 36538 39488 36544 39500
rect 35912 39460 36544 39488
rect 33781 39451 33839 39457
rect 36538 39448 36544 39460
rect 36596 39448 36602 39500
rect 36722 39448 36728 39500
rect 36780 39448 36786 39500
rect 38102 39448 38108 39500
rect 38160 39488 38166 39500
rect 40052 39488 40080 39596
rect 40954 39516 40960 39568
rect 41012 39556 41018 39568
rect 41064 39556 41092 39596
rect 41432 39596 42901 39624
rect 41432 39565 41460 39596
rect 42889 39593 42901 39596
rect 42935 39593 42947 39627
rect 42889 39587 42947 39593
rect 42978 39584 42984 39636
rect 43036 39624 43042 39636
rect 43717 39627 43775 39633
rect 43717 39624 43729 39627
rect 43036 39596 43729 39624
rect 43036 39584 43042 39596
rect 43717 39593 43729 39596
rect 43763 39593 43775 39627
rect 43717 39587 43775 39593
rect 44082 39584 44088 39636
rect 44140 39624 44146 39636
rect 44177 39627 44235 39633
rect 44177 39624 44189 39627
rect 44140 39596 44189 39624
rect 44140 39584 44146 39596
rect 44177 39593 44189 39596
rect 44223 39593 44235 39627
rect 44177 39587 44235 39593
rect 46106 39584 46112 39636
rect 46164 39584 46170 39636
rect 46477 39627 46535 39633
rect 46477 39593 46489 39627
rect 46523 39624 46535 39627
rect 46658 39624 46664 39636
rect 46523 39596 46664 39624
rect 46523 39593 46535 39596
rect 46477 39587 46535 39593
rect 46658 39584 46664 39596
rect 46716 39584 46722 39636
rect 48406 39584 48412 39636
rect 48464 39624 48470 39636
rect 49878 39624 49884 39636
rect 48464 39596 49884 39624
rect 48464 39584 48470 39596
rect 49878 39584 49884 39596
rect 49936 39584 49942 39636
rect 49970 39584 49976 39636
rect 50028 39624 50034 39636
rect 50028 39596 51074 39624
rect 50028 39584 50034 39596
rect 41012 39528 41092 39556
rect 41417 39559 41475 39565
rect 41012 39516 41018 39528
rect 41417 39525 41429 39559
rect 41463 39525 41475 39559
rect 41417 39519 41475 39525
rect 41506 39516 41512 39568
rect 41564 39556 41570 39568
rect 43257 39559 43315 39565
rect 43257 39556 43269 39559
rect 41564 39528 43269 39556
rect 41564 39516 41570 39528
rect 43257 39525 43269 39528
rect 43303 39525 43315 39559
rect 43257 39519 43315 39525
rect 43438 39516 43444 39568
rect 43496 39556 43502 39568
rect 45738 39556 45744 39568
rect 43496 39528 45744 39556
rect 43496 39516 43502 39528
rect 45738 39516 45744 39528
rect 45796 39556 45802 39568
rect 45796 39528 45968 39556
rect 45796 39516 45802 39528
rect 38160 39460 40080 39488
rect 41693 39491 41751 39497
rect 38160 39448 38166 39460
rect 41693 39457 41705 39491
rect 41739 39488 41751 39491
rect 41739 39460 41828 39488
rect 41739 39457 41751 39460
rect 41693 39451 41751 39457
rect 41800 39432 41828 39460
rect 42426 39448 42432 39500
rect 42484 39448 42490 39500
rect 42521 39491 42579 39497
rect 42521 39457 42533 39491
rect 42567 39488 42579 39491
rect 42702 39488 42708 39500
rect 42567 39460 42708 39488
rect 42567 39457 42579 39460
rect 42521 39451 42579 39457
rect 42702 39448 42708 39460
rect 42760 39448 42766 39500
rect 44085 39491 44143 39497
rect 43272 39460 43576 39488
rect 30098 39380 30104 39432
rect 30156 39420 30162 39432
rect 30745 39423 30803 39429
rect 30745 39420 30757 39423
rect 30156 39392 30757 39420
rect 30156 39380 30162 39392
rect 30745 39389 30757 39392
rect 30791 39420 30803 39423
rect 30834 39420 30840 39432
rect 30791 39392 30840 39420
rect 30791 39389 30803 39392
rect 30745 39383 30803 39389
rect 30834 39380 30840 39392
rect 30892 39380 30898 39432
rect 30929 39423 30987 39429
rect 30929 39389 30941 39423
rect 30975 39389 30987 39423
rect 31849 39423 31907 39429
rect 31849 39420 31861 39423
rect 30929 39383 30987 39389
rect 31404 39392 31861 39420
rect 27948 39324 30052 39352
rect 27948 39312 27954 39324
rect 20588 39256 22094 39284
rect 20588 39244 20594 39256
rect 24118 39244 24124 39296
rect 24176 39284 24182 39296
rect 24397 39287 24455 39293
rect 24397 39284 24409 39287
rect 24176 39256 24409 39284
rect 24176 39244 24182 39256
rect 24397 39253 24409 39256
rect 24443 39253 24455 39287
rect 24397 39247 24455 39253
rect 25958 39244 25964 39296
rect 26016 39284 26022 39296
rect 26421 39287 26479 39293
rect 26421 39284 26433 39287
rect 26016 39256 26433 39284
rect 26016 39244 26022 39256
rect 26421 39253 26433 39256
rect 26467 39253 26479 39287
rect 26421 39247 26479 39253
rect 26510 39244 26516 39296
rect 26568 39284 26574 39296
rect 27157 39287 27215 39293
rect 27157 39284 27169 39287
rect 26568 39256 27169 39284
rect 26568 39244 26574 39256
rect 27157 39253 27169 39256
rect 27203 39253 27215 39287
rect 27157 39247 27215 39253
rect 27246 39244 27252 39296
rect 27304 39284 27310 39296
rect 28994 39284 29000 39296
rect 27304 39256 29000 39284
rect 27304 39244 27310 39256
rect 28994 39244 29000 39256
rect 29052 39244 29058 39296
rect 29086 39244 29092 39296
rect 29144 39284 29150 39296
rect 29273 39287 29331 39293
rect 29273 39284 29285 39287
rect 29144 39256 29285 39284
rect 29144 39244 29150 39256
rect 29273 39253 29285 39256
rect 29319 39253 29331 39287
rect 30944 39284 30972 39383
rect 31404 39361 31432 39392
rect 31849 39389 31861 39392
rect 31895 39389 31907 39423
rect 31849 39383 31907 39389
rect 32214 39380 32220 39432
rect 32272 39420 32278 39432
rect 32582 39420 32588 39432
rect 32272 39392 32588 39420
rect 32272 39380 32278 39392
rect 32582 39380 32588 39392
rect 32640 39420 32646 39432
rect 33965 39423 34023 39429
rect 33965 39420 33977 39423
rect 32640 39392 33977 39420
rect 32640 39380 32646 39392
rect 33965 39389 33977 39392
rect 34011 39420 34023 39423
rect 35897 39423 35955 39429
rect 35897 39420 35909 39423
rect 34011 39392 35909 39420
rect 34011 39389 34023 39392
rect 33965 39383 34023 39389
rect 35897 39389 35909 39392
rect 35943 39420 35955 39423
rect 37366 39420 37372 39432
rect 35943 39392 37372 39420
rect 35943 39389 35955 39392
rect 35897 39383 35955 39389
rect 37366 39380 37372 39392
rect 37424 39380 37430 39432
rect 37458 39380 37464 39432
rect 37516 39420 37522 39432
rect 38562 39420 38568 39432
rect 37516 39392 38568 39420
rect 37516 39380 37522 39392
rect 38562 39380 38568 39392
rect 38620 39380 38626 39432
rect 39114 39380 39120 39432
rect 39172 39380 39178 39432
rect 41414 39420 41420 39432
rect 39960 39392 41420 39420
rect 31389 39355 31447 39361
rect 31389 39321 31401 39355
rect 31435 39321 31447 39355
rect 31389 39315 31447 39321
rect 33226 39312 33232 39364
rect 33284 39352 33290 39364
rect 33284 39324 35572 39352
rect 33284 39312 33290 39324
rect 32398 39284 32404 39296
rect 30944 39256 32404 39284
rect 29273 39247 29331 39253
rect 32398 39244 32404 39256
rect 32456 39244 32462 39296
rect 33321 39287 33379 39293
rect 33321 39253 33333 39287
rect 33367 39284 33379 39287
rect 33502 39284 33508 39296
rect 33367 39256 33508 39284
rect 33367 39253 33379 39256
rect 33321 39247 33379 39253
rect 33502 39244 33508 39256
rect 33560 39244 33566 39296
rect 35544 39284 35572 39324
rect 35618 39312 35624 39364
rect 35676 39352 35682 39364
rect 36722 39352 36728 39364
rect 35676 39324 36728 39352
rect 35676 39312 35682 39324
rect 36722 39312 36728 39324
rect 36780 39312 36786 39364
rect 39960 39361 39988 39392
rect 41414 39380 41420 39392
rect 41472 39380 41478 39432
rect 41782 39380 41788 39432
rect 41840 39380 41846 39432
rect 41874 39380 41880 39432
rect 41932 39420 41938 39432
rect 42610 39420 42616 39432
rect 41932 39392 42616 39420
rect 41932 39380 41938 39392
rect 42610 39380 42616 39392
rect 42668 39420 42674 39432
rect 43272 39420 43300 39460
rect 42668 39392 43300 39420
rect 43349 39423 43407 39429
rect 42668 39380 42674 39392
rect 43349 39389 43361 39423
rect 43395 39389 43407 39423
rect 43349 39383 43407 39389
rect 39945 39355 40003 39361
rect 39945 39352 39957 39355
rect 38028 39324 39957 39352
rect 37458 39284 37464 39296
rect 35544 39256 37464 39284
rect 37458 39244 37464 39256
rect 37516 39244 37522 39296
rect 37550 39244 37556 39296
rect 37608 39284 37614 39296
rect 38028 39284 38056 39324
rect 39945 39321 39957 39324
rect 39991 39321 40003 39355
rect 40402 39352 40408 39364
rect 39945 39315 40003 39321
rect 40052 39324 40408 39352
rect 37608 39256 38056 39284
rect 38473 39287 38531 39293
rect 37608 39244 37614 39256
rect 38473 39253 38485 39287
rect 38519 39284 38531 39287
rect 38746 39284 38752 39296
rect 38519 39256 38752 39284
rect 38519 39253 38531 39256
rect 38473 39247 38531 39253
rect 38746 39244 38752 39256
rect 38804 39284 38810 39296
rect 40052 39284 40080 39324
rect 40402 39312 40408 39324
rect 40460 39312 40466 39364
rect 41966 39352 41972 39364
rect 41708 39324 41972 39352
rect 38804 39256 40080 39284
rect 38804 39244 38810 39256
rect 40126 39244 40132 39296
rect 40184 39284 40190 39296
rect 41046 39284 41052 39296
rect 40184 39256 41052 39284
rect 40184 39244 40190 39256
rect 41046 39244 41052 39256
rect 41104 39284 41110 39296
rect 41708 39284 41736 39324
rect 41966 39312 41972 39324
rect 42024 39312 42030 39364
rect 42150 39312 42156 39364
rect 42208 39352 42214 39364
rect 43364 39352 43392 39383
rect 43438 39380 43444 39432
rect 43496 39380 43502 39432
rect 43548 39420 43576 39460
rect 44085 39457 44097 39491
rect 44131 39488 44143 39491
rect 45278 39488 45284 39500
rect 44131 39460 45284 39488
rect 44131 39457 44143 39460
rect 44085 39451 44143 39457
rect 45278 39448 45284 39460
rect 45336 39448 45342 39500
rect 45649 39491 45707 39497
rect 45649 39488 45661 39491
rect 45388 39460 45661 39488
rect 44269 39423 44327 39429
rect 44269 39420 44281 39423
rect 43548 39392 44281 39420
rect 44269 39389 44281 39392
rect 44315 39389 44327 39423
rect 44269 39383 44327 39389
rect 45094 39380 45100 39432
rect 45152 39420 45158 39432
rect 45388 39420 45416 39460
rect 45649 39457 45661 39460
rect 45695 39488 45707 39491
rect 45830 39488 45836 39500
rect 45695 39460 45836 39488
rect 45695 39457 45707 39460
rect 45649 39451 45707 39457
rect 45830 39448 45836 39460
rect 45888 39448 45894 39500
rect 45940 39488 45968 39528
rect 46014 39516 46020 39568
rect 46072 39556 46078 39568
rect 46072 39528 47072 39556
rect 46072 39516 46078 39528
rect 46290 39488 46296 39500
rect 45940 39460 46296 39488
rect 46290 39448 46296 39460
rect 46348 39448 46354 39500
rect 47044 39497 47072 39528
rect 48314 39516 48320 39568
rect 48372 39556 48378 39568
rect 48866 39556 48872 39568
rect 48372 39528 48872 39556
rect 48372 39516 48378 39528
rect 48866 39516 48872 39528
rect 48924 39556 48930 39568
rect 48924 39528 49082 39556
rect 48924 39516 48930 39528
rect 50246 39516 50252 39568
rect 50304 39516 50310 39568
rect 50614 39516 50620 39568
rect 50672 39516 50678 39568
rect 47029 39491 47087 39497
rect 47029 39457 47041 39491
rect 47075 39488 47087 39491
rect 48774 39488 48780 39500
rect 47075 39460 48780 39488
rect 47075 39457 47087 39460
rect 47029 39451 47087 39457
rect 48774 39448 48780 39460
rect 48832 39448 48838 39500
rect 51046 39488 51074 39596
rect 52362 39584 52368 39636
rect 52420 39584 52426 39636
rect 52730 39584 52736 39636
rect 52788 39624 52794 39636
rect 63494 39624 63500 39636
rect 52788 39596 63500 39624
rect 52788 39584 52794 39596
rect 63494 39584 63500 39596
rect 63552 39584 63558 39636
rect 51350 39516 51356 39568
rect 51408 39556 51414 39568
rect 52178 39556 52184 39568
rect 51408 39528 52184 39556
rect 51408 39516 51414 39528
rect 52178 39516 52184 39528
rect 52236 39516 52242 39568
rect 52822 39516 52828 39568
rect 52880 39516 52886 39568
rect 54754 39516 54760 39568
rect 54812 39556 54818 39568
rect 54812 39528 58572 39556
rect 54812 39516 54818 39528
rect 51169 39491 51227 39497
rect 51169 39488 51181 39491
rect 51046 39460 51181 39488
rect 51169 39457 51181 39460
rect 51215 39457 51227 39491
rect 51169 39451 51227 39457
rect 52086 39448 52092 39500
rect 52144 39488 52150 39500
rect 52638 39488 52644 39500
rect 52144 39460 52644 39488
rect 52144 39448 52150 39460
rect 52638 39448 52644 39460
rect 52696 39488 52702 39500
rect 52733 39491 52791 39497
rect 52733 39488 52745 39491
rect 52696 39460 52745 39488
rect 52696 39448 52702 39460
rect 52733 39457 52745 39460
rect 52779 39457 52791 39491
rect 54662 39488 54668 39500
rect 52733 39451 52791 39457
rect 53024 39460 54668 39488
rect 45152 39392 45416 39420
rect 45465 39423 45523 39429
rect 45152 39380 45158 39392
rect 45465 39389 45477 39423
rect 45511 39389 45523 39423
rect 45465 39383 45523 39389
rect 42208 39324 43392 39352
rect 45480 39352 45508 39383
rect 45554 39380 45560 39432
rect 45612 39380 45618 39432
rect 46569 39423 46627 39429
rect 46569 39420 46581 39423
rect 46032 39392 46581 39420
rect 45922 39352 45928 39364
rect 45480 39324 45928 39352
rect 42208 39312 42214 39324
rect 45922 39312 45928 39324
rect 45980 39312 45986 39364
rect 46032 39361 46060 39392
rect 46569 39389 46581 39392
rect 46615 39389 46627 39423
rect 46569 39383 46627 39389
rect 46750 39380 46756 39432
rect 46808 39380 46814 39432
rect 48406 39420 48412 39432
rect 47320 39392 48412 39420
rect 46017 39355 46075 39361
rect 46017 39321 46029 39355
rect 46063 39321 46075 39355
rect 46017 39315 46075 39321
rect 41104 39256 41736 39284
rect 41104 39244 41110 39256
rect 41782 39244 41788 39296
rect 41840 39284 41846 39296
rect 42061 39287 42119 39293
rect 42061 39284 42073 39287
rect 41840 39256 42073 39284
rect 41840 39244 41846 39256
rect 42061 39253 42073 39256
rect 42107 39253 42119 39287
rect 42061 39247 42119 39253
rect 42334 39244 42340 39296
rect 42392 39284 42398 39296
rect 47320 39284 47348 39392
rect 48406 39380 48412 39392
rect 48464 39420 48470 39432
rect 48501 39423 48559 39429
rect 48501 39420 48513 39423
rect 48464 39392 48513 39420
rect 48464 39380 48470 39392
rect 48501 39389 48513 39392
rect 48547 39389 48559 39423
rect 50525 39423 50583 39429
rect 50525 39420 50537 39423
rect 48501 39383 48559 39389
rect 48792 39392 50537 39420
rect 48130 39312 48136 39364
rect 48188 39352 48194 39364
rect 48792 39352 48820 39392
rect 50525 39389 50537 39392
rect 50571 39420 50583 39423
rect 50706 39420 50712 39432
rect 50571 39392 50712 39420
rect 50571 39389 50583 39392
rect 50525 39383 50583 39389
rect 50706 39380 50712 39392
rect 50764 39380 50770 39432
rect 53024 39429 53052 39460
rect 54662 39448 54668 39460
rect 54720 39448 54726 39500
rect 58544 39497 58572 39528
rect 59262 39516 59268 39568
rect 59320 39516 59326 39568
rect 55861 39491 55919 39497
rect 55861 39457 55873 39491
rect 55907 39488 55919 39491
rect 56413 39491 56471 39497
rect 56413 39488 56425 39491
rect 55907 39460 56425 39488
rect 55907 39457 55919 39460
rect 55861 39451 55919 39457
rect 56413 39457 56425 39460
rect 56459 39457 56471 39491
rect 56413 39451 56471 39457
rect 58529 39491 58587 39497
rect 58529 39457 58541 39491
rect 58575 39457 58587 39491
rect 58529 39451 58587 39457
rect 53009 39423 53067 39429
rect 53009 39389 53021 39423
rect 53055 39389 53067 39423
rect 53009 39383 53067 39389
rect 53558 39380 53564 39432
rect 53616 39420 53622 39432
rect 53837 39423 53895 39429
rect 53837 39420 53849 39423
rect 53616 39392 53849 39420
rect 53616 39380 53622 39392
rect 53837 39389 53849 39392
rect 53883 39389 53895 39423
rect 53837 39383 53895 39389
rect 55950 39380 55956 39432
rect 56008 39380 56014 39432
rect 56137 39423 56195 39429
rect 56137 39389 56149 39423
rect 56183 39420 56195 39423
rect 56318 39420 56324 39432
rect 56183 39392 56324 39420
rect 56183 39389 56195 39392
rect 56137 39383 56195 39389
rect 56318 39380 56324 39392
rect 56376 39380 56382 39432
rect 56778 39380 56784 39432
rect 56836 39420 56842 39432
rect 56965 39423 57023 39429
rect 56965 39420 56977 39423
rect 56836 39392 56977 39420
rect 56836 39380 56842 39392
rect 56965 39389 56977 39392
rect 57011 39389 57023 39423
rect 56965 39383 57023 39389
rect 58805 39423 58863 39429
rect 58805 39389 58817 39423
rect 58851 39420 58863 39423
rect 60921 39423 60979 39429
rect 60921 39420 60933 39423
rect 58851 39392 59952 39420
rect 58851 39389 58863 39392
rect 58805 39383 58863 39389
rect 59924 39364 59952 39392
rect 60292 39392 60933 39420
rect 48188 39324 48820 39352
rect 48188 39312 48194 39324
rect 50798 39312 50804 39364
rect 50856 39352 50862 39364
rect 56686 39352 56692 39364
rect 50856 39324 56692 39352
rect 50856 39312 50862 39324
rect 56686 39312 56692 39324
rect 56744 39312 56750 39364
rect 59906 39312 59912 39364
rect 59964 39312 59970 39364
rect 60292 39296 60320 39392
rect 60921 39389 60933 39392
rect 60967 39389 60979 39423
rect 60921 39383 60979 39389
rect 42392 39256 47348 39284
rect 42392 39244 42398 39256
rect 47394 39244 47400 39296
rect 47452 39284 47458 39296
rect 47673 39287 47731 39293
rect 47673 39284 47685 39287
rect 47452 39256 47685 39284
rect 47452 39244 47458 39256
rect 47673 39253 47685 39256
rect 47719 39253 47731 39287
rect 47673 39247 47731 39253
rect 53190 39244 53196 39296
rect 53248 39244 53254 39296
rect 55306 39244 55312 39296
rect 55364 39284 55370 39296
rect 55493 39287 55551 39293
rect 55493 39284 55505 39287
rect 55364 39256 55505 39284
rect 55364 39244 55370 39256
rect 55493 39253 55505 39256
rect 55539 39253 55551 39287
rect 55493 39247 55551 39253
rect 56226 39244 56232 39296
rect 56284 39284 56290 39296
rect 59170 39284 59176 39296
rect 56284 39256 59176 39284
rect 56284 39244 56290 39256
rect 59170 39244 59176 39256
rect 59228 39244 59234 39296
rect 60274 39244 60280 39296
rect 60332 39244 60338 39296
rect 60366 39244 60372 39296
rect 60424 39244 60430 39296
rect 552 39194 66424 39216
rect 552 39142 1998 39194
rect 2050 39142 2062 39194
rect 2114 39142 2126 39194
rect 2178 39142 2190 39194
rect 2242 39142 2254 39194
rect 2306 39142 49998 39194
rect 50050 39142 50062 39194
rect 50114 39142 50126 39194
rect 50178 39142 50190 39194
rect 50242 39142 50254 39194
rect 50306 39142 66424 39194
rect 552 39120 66424 39142
rect 8570 39040 8576 39092
rect 8628 39080 8634 39092
rect 11422 39080 11428 39092
rect 8628 39052 9996 39080
rect 8628 39040 8634 39052
rect 8481 38947 8539 38953
rect 8481 38913 8493 38947
rect 8527 38944 8539 38947
rect 8754 38944 8760 38956
rect 8527 38916 8760 38944
rect 8527 38913 8539 38916
rect 8481 38907 8539 38913
rect 8754 38904 8760 38916
rect 8812 38904 8818 38956
rect 8205 38879 8263 38885
rect 8205 38845 8217 38879
rect 8251 38845 8263 38879
rect 8205 38839 8263 38845
rect 8220 38808 8248 38839
rect 8662 38808 8668 38820
rect 8220 38780 8668 38808
rect 8662 38768 8668 38780
rect 8720 38768 8726 38820
rect 8757 38811 8815 38817
rect 8757 38777 8769 38811
rect 8803 38808 8815 38811
rect 8846 38808 8852 38820
rect 8803 38780 8852 38808
rect 8803 38777 8815 38780
rect 8757 38771 8815 38777
rect 8846 38768 8852 38780
rect 8904 38768 8910 38820
rect 9968 38808 9996 39052
rect 10520 39052 11428 39080
rect 10520 38953 10548 39052
rect 11422 39040 11428 39052
rect 11480 39040 11486 39092
rect 12912 39052 15240 39080
rect 10505 38947 10563 38953
rect 10505 38913 10517 38947
rect 10551 38913 10563 38947
rect 10505 38907 10563 38913
rect 10597 38947 10655 38953
rect 10597 38913 10609 38947
rect 10643 38944 10655 38947
rect 11514 38944 11520 38956
rect 10643 38916 11520 38944
rect 10643 38913 10655 38916
rect 10597 38907 10655 38913
rect 11514 38904 11520 38916
rect 11572 38944 11578 38956
rect 11572 38916 12204 38944
rect 11572 38904 11578 38916
rect 9968 38794 10548 38808
rect 9982 38780 10548 38794
rect 7558 38700 7564 38752
rect 7616 38700 7622 38752
rect 10520 38740 10548 38780
rect 10870 38768 10876 38820
rect 10928 38768 10934 38820
rect 10962 38768 10968 38820
rect 11020 38808 11026 38820
rect 12176 38808 12204 38916
rect 12802 38904 12808 38956
rect 12860 38904 12866 38956
rect 12912 38953 12940 39052
rect 15212 39024 15240 39052
rect 20162 39040 20168 39092
rect 20220 39080 20226 39092
rect 21177 39083 21235 39089
rect 21177 39080 21189 39083
rect 20220 39052 21189 39080
rect 20220 39040 20226 39052
rect 21177 39049 21189 39052
rect 21223 39049 21235 39083
rect 21177 39043 21235 39049
rect 23661 39083 23719 39089
rect 23661 39049 23673 39083
rect 23707 39080 23719 39083
rect 23934 39080 23940 39092
rect 23707 39052 23940 39080
rect 23707 39049 23719 39052
rect 23661 39043 23719 39049
rect 23934 39040 23940 39052
rect 23992 39040 23998 39092
rect 24302 39040 24308 39092
rect 24360 39080 24366 39092
rect 24360 39052 25636 39080
rect 24360 39040 24366 39052
rect 25608 39024 25636 39052
rect 26050 39040 26056 39092
rect 26108 39080 26114 39092
rect 26108 39052 27752 39080
rect 26108 39040 26114 39052
rect 15194 38972 15200 39024
rect 15252 39012 15258 39024
rect 15289 39015 15347 39021
rect 15289 39012 15301 39015
rect 15252 38984 15301 39012
rect 15252 38972 15258 38984
rect 15289 38981 15301 38984
rect 15335 39012 15347 39015
rect 16390 39012 16396 39024
rect 15335 38984 16396 39012
rect 15335 38981 15347 38984
rect 15289 38975 15347 38981
rect 16390 38972 16396 38984
rect 16448 38972 16454 39024
rect 21085 39015 21143 39021
rect 21085 38981 21097 39015
rect 21131 39012 21143 39015
rect 21726 39012 21732 39024
rect 21131 38984 21732 39012
rect 21131 38981 21143 38984
rect 21085 38975 21143 38981
rect 21726 38972 21732 38984
rect 21784 38972 21790 39024
rect 25590 38972 25596 39024
rect 25648 39012 25654 39024
rect 26694 39012 26700 39024
rect 25648 38984 26700 39012
rect 25648 38972 25654 38984
rect 26694 38972 26700 38984
rect 26752 38972 26758 39024
rect 12897 38947 12955 38953
rect 12897 38913 12909 38947
rect 12943 38913 12955 38947
rect 12897 38907 12955 38913
rect 13541 38947 13599 38953
rect 13541 38913 13553 38947
rect 13587 38944 13599 38947
rect 13814 38944 13820 38956
rect 13587 38916 13820 38944
rect 13587 38913 13599 38916
rect 13541 38907 13599 38913
rect 13814 38904 13820 38916
rect 13872 38944 13878 38956
rect 14826 38944 14832 38956
rect 13872 38916 14832 38944
rect 13872 38904 13878 38916
rect 14826 38904 14832 38916
rect 14884 38944 14890 38956
rect 16758 38944 16764 38956
rect 14884 38916 16764 38944
rect 14884 38904 14890 38916
rect 16758 38904 16764 38916
rect 16816 38904 16822 38956
rect 19058 38904 19064 38956
rect 19116 38944 19122 38956
rect 19337 38947 19395 38953
rect 19337 38944 19349 38947
rect 19116 38916 19349 38944
rect 19116 38904 19122 38916
rect 19337 38913 19349 38916
rect 19383 38944 19395 38947
rect 21910 38944 21916 38956
rect 19383 38916 21916 38944
rect 19383 38913 19395 38916
rect 19337 38907 19395 38913
rect 21910 38904 21916 38916
rect 21968 38904 21974 38956
rect 22186 38904 22192 38956
rect 22244 38944 22250 38956
rect 23382 38944 23388 38956
rect 22244 38916 23388 38944
rect 22244 38904 22250 38916
rect 23382 38904 23388 38916
rect 23440 38944 23446 38956
rect 23845 38947 23903 38953
rect 23845 38944 23857 38947
rect 23440 38916 23857 38944
rect 23440 38904 23446 38916
rect 23845 38913 23857 38916
rect 23891 38913 23903 38947
rect 23845 38907 23903 38913
rect 24118 38904 24124 38956
rect 24176 38904 24182 38956
rect 24210 38904 24216 38956
rect 24268 38944 24274 38956
rect 24486 38944 24492 38956
rect 24268 38916 24492 38944
rect 24268 38904 24274 38916
rect 24486 38904 24492 38916
rect 24544 38944 24550 38956
rect 26329 38947 26387 38953
rect 26329 38944 26341 38947
rect 24544 38916 26341 38944
rect 24544 38904 24550 38916
rect 26329 38913 26341 38916
rect 26375 38944 26387 38947
rect 27617 38947 27675 38953
rect 27617 38944 27629 38947
rect 26375 38916 27629 38944
rect 26375 38913 26387 38916
rect 26329 38907 26387 38913
rect 27617 38913 27629 38916
rect 27663 38913 27675 38947
rect 27724 38944 27752 39052
rect 27982 39040 27988 39092
rect 28040 39080 28046 39092
rect 42334 39080 42340 39092
rect 28040 39052 42340 39080
rect 28040 39040 28046 39052
rect 42334 39040 42340 39052
rect 42392 39040 42398 39092
rect 42426 39040 42432 39092
rect 42484 39080 42490 39092
rect 43349 39083 43407 39089
rect 43349 39080 43361 39083
rect 42484 39052 43361 39080
rect 42484 39040 42490 39052
rect 43349 39049 43361 39052
rect 43395 39049 43407 39083
rect 43349 39043 43407 39049
rect 45278 39040 45284 39092
rect 45336 39040 45342 39092
rect 46014 39040 46020 39092
rect 46072 39080 46078 39092
rect 46109 39083 46167 39089
rect 46109 39080 46121 39083
rect 46072 39052 46121 39080
rect 46072 39040 46078 39052
rect 46109 39049 46121 39052
rect 46155 39049 46167 39083
rect 46109 39043 46167 39049
rect 48685 39083 48743 39089
rect 48685 39049 48697 39083
rect 48731 39080 48743 39083
rect 49050 39080 49056 39092
rect 48731 39052 49056 39080
rect 48731 39049 48743 39052
rect 48685 39043 48743 39049
rect 49050 39040 49056 39052
rect 49108 39040 49114 39092
rect 60458 39080 60464 39092
rect 58636 39052 60464 39080
rect 28000 38984 28580 39012
rect 28000 38944 28028 38984
rect 28552 38953 28580 38984
rect 30392 38984 31064 39012
rect 27724 38916 28028 38944
rect 28537 38947 28595 38953
rect 27617 38907 27675 38913
rect 28537 38913 28549 38947
rect 28583 38944 28595 38947
rect 30098 38944 30104 38956
rect 28583 38916 30104 38944
rect 28583 38913 28595 38916
rect 28537 38907 28595 38913
rect 30098 38904 30104 38916
rect 30156 38904 30162 38956
rect 30193 38947 30251 38953
rect 30193 38913 30205 38947
rect 30239 38944 30251 38947
rect 30282 38944 30288 38956
rect 30239 38916 30288 38944
rect 30239 38913 30251 38916
rect 30193 38907 30251 38913
rect 30282 38904 30288 38916
rect 30340 38904 30346 38956
rect 12986 38836 12992 38888
rect 13044 38836 13050 38888
rect 15286 38836 15292 38888
rect 15344 38876 15350 38888
rect 16025 38879 16083 38885
rect 16025 38876 16037 38879
rect 15344 38848 16037 38876
rect 15344 38836 15350 38848
rect 16025 38845 16037 38848
rect 16071 38845 16083 38879
rect 16025 38839 16083 38845
rect 21726 38836 21732 38888
rect 21784 38836 21790 38888
rect 26053 38879 26111 38885
rect 26053 38845 26065 38879
rect 26099 38876 26111 38879
rect 26510 38876 26516 38888
rect 26099 38848 26516 38876
rect 26099 38845 26111 38848
rect 26053 38839 26111 38845
rect 26510 38836 26516 38848
rect 26568 38836 26574 38888
rect 26694 38836 26700 38888
rect 26752 38876 26758 38888
rect 30392 38876 30420 38984
rect 30466 38904 30472 38956
rect 30524 38944 30530 38956
rect 30929 38947 30987 38953
rect 30929 38944 30941 38947
rect 30524 38916 30941 38944
rect 30524 38904 30530 38916
rect 30929 38913 30941 38916
rect 30975 38913 30987 38947
rect 31036 38944 31064 38984
rect 31110 38972 31116 39024
rect 31168 39012 31174 39024
rect 31573 39015 31631 39021
rect 31573 39012 31585 39015
rect 31168 38984 31585 39012
rect 31168 38972 31174 38984
rect 31573 38981 31585 38984
rect 31619 38981 31631 39015
rect 33594 39012 33600 39024
rect 31573 38975 31631 38981
rect 31680 38984 33600 39012
rect 31680 38944 31708 38984
rect 33594 38972 33600 38984
rect 33652 38972 33658 39024
rect 37550 39012 37556 39024
rect 34256 38984 35756 39012
rect 31036 38916 31708 38944
rect 30929 38907 30987 38913
rect 32214 38904 32220 38956
rect 32272 38904 32278 38956
rect 26752 38848 30420 38876
rect 30745 38879 30803 38885
rect 26752 38836 26758 38848
rect 30745 38845 30757 38879
rect 30791 38876 30803 38879
rect 31662 38876 31668 38888
rect 30791 38848 31668 38876
rect 30791 38845 30803 38848
rect 30745 38839 30803 38845
rect 31662 38836 31668 38848
rect 31720 38876 31726 38888
rect 32033 38879 32091 38885
rect 32033 38876 32045 38879
rect 31720 38848 32045 38876
rect 31720 38836 31726 38848
rect 32033 38845 32045 38848
rect 32079 38845 32091 38879
rect 32033 38839 32091 38845
rect 32398 38836 32404 38888
rect 32456 38836 32462 38888
rect 32953 38879 33011 38885
rect 32953 38845 32965 38879
rect 32999 38876 33011 38879
rect 32999 38848 33548 38876
rect 32999 38845 33011 38848
rect 32953 38839 33011 38845
rect 13446 38808 13452 38820
rect 11020 38780 11362 38808
rect 12176 38780 13452 38808
rect 11020 38768 11026 38780
rect 13446 38768 13452 38780
rect 13504 38768 13510 38820
rect 13817 38811 13875 38817
rect 13817 38777 13829 38811
rect 13863 38777 13875 38811
rect 13817 38771 13875 38777
rect 10980 38740 11008 38768
rect 10520 38712 11008 38740
rect 12342 38700 12348 38752
rect 12400 38700 12406 38752
rect 13357 38743 13415 38749
rect 13357 38709 13369 38743
rect 13403 38740 13415 38743
rect 13832 38740 13860 38771
rect 14090 38768 14096 38820
rect 14148 38808 14154 38820
rect 18509 38811 18567 38817
rect 14148 38780 14306 38808
rect 14148 38768 14154 38780
rect 18509 38777 18521 38811
rect 18555 38808 18567 38811
rect 19518 38808 19524 38820
rect 18555 38780 19524 38808
rect 18555 38777 18567 38780
rect 18509 38771 18567 38777
rect 19518 38768 19524 38780
rect 19576 38768 19582 38820
rect 19610 38768 19616 38820
rect 19668 38768 19674 38820
rect 19720 38780 20102 38808
rect 13403 38712 13860 38740
rect 13403 38709 13415 38712
rect 13357 38703 13415 38709
rect 15378 38700 15384 38752
rect 15436 38740 15442 38752
rect 15473 38743 15531 38749
rect 15473 38740 15485 38743
rect 15436 38712 15485 38740
rect 15436 38700 15442 38712
rect 15473 38709 15485 38712
rect 15519 38709 15531 38743
rect 15473 38703 15531 38709
rect 18046 38700 18052 38752
rect 18104 38740 18110 38752
rect 19242 38740 19248 38752
rect 18104 38712 19248 38740
rect 18104 38700 18110 38712
rect 19242 38700 19248 38712
rect 19300 38740 19306 38752
rect 19720 38740 19748 38780
rect 19300 38712 19748 38740
rect 19996 38740 20024 38780
rect 22186 38768 22192 38820
rect 22244 38768 22250 38820
rect 27433 38811 27491 38817
rect 23414 38780 24610 38808
rect 21358 38740 21364 38752
rect 19996 38712 21364 38740
rect 19300 38700 19306 38712
rect 21358 38700 21364 38712
rect 21416 38740 21422 38752
rect 22002 38740 22008 38752
rect 21416 38712 22008 38740
rect 21416 38700 21422 38712
rect 22002 38700 22008 38712
rect 22060 38700 22066 38752
rect 24504 38740 24532 38780
rect 27433 38777 27445 38811
rect 27479 38808 27491 38811
rect 28902 38808 28908 38820
rect 27479 38780 28908 38808
rect 27479 38777 27491 38780
rect 27433 38771 27491 38777
rect 28902 38768 28908 38780
rect 28960 38768 28966 38820
rect 28994 38768 29000 38820
rect 29052 38808 29058 38820
rect 29052 38780 30512 38808
rect 29052 38768 29058 38780
rect 24946 38740 24952 38752
rect 24504 38712 24952 38740
rect 24946 38700 24952 38712
rect 25004 38700 25010 38752
rect 25682 38700 25688 38752
rect 25740 38700 25746 38752
rect 26142 38700 26148 38752
rect 26200 38700 26206 38752
rect 26786 38700 26792 38752
rect 26844 38740 26850 38752
rect 27065 38743 27123 38749
rect 27065 38740 27077 38743
rect 26844 38712 27077 38740
rect 26844 38700 26850 38712
rect 27065 38709 27077 38712
rect 27111 38709 27123 38743
rect 27065 38703 27123 38709
rect 27525 38743 27583 38749
rect 27525 38709 27537 38743
rect 27571 38740 27583 38743
rect 27706 38740 27712 38752
rect 27571 38712 27712 38740
rect 27571 38709 27583 38712
rect 27525 38703 27583 38709
rect 27706 38700 27712 38712
rect 27764 38700 27770 38752
rect 27798 38700 27804 38752
rect 27856 38740 27862 38752
rect 27893 38743 27951 38749
rect 27893 38740 27905 38743
rect 27856 38712 27905 38740
rect 27856 38700 27862 38712
rect 27893 38709 27905 38712
rect 27939 38709 27951 38743
rect 27893 38703 27951 38709
rect 28258 38700 28264 38752
rect 28316 38700 28322 38752
rect 28353 38743 28411 38749
rect 28353 38709 28365 38743
rect 28399 38740 28411 38743
rect 29086 38740 29092 38752
rect 28399 38712 29092 38740
rect 28399 38709 28411 38712
rect 28353 38703 28411 38709
rect 29086 38700 29092 38712
rect 29144 38700 29150 38752
rect 29178 38700 29184 38752
rect 29236 38740 29242 38752
rect 29549 38743 29607 38749
rect 29549 38740 29561 38743
rect 29236 38712 29561 38740
rect 29236 38700 29242 38712
rect 29549 38709 29561 38712
rect 29595 38709 29607 38743
rect 29549 38703 29607 38709
rect 29914 38700 29920 38752
rect 29972 38700 29978 38752
rect 30009 38743 30067 38749
rect 30009 38709 30021 38743
rect 30055 38740 30067 38743
rect 30377 38743 30435 38749
rect 30377 38740 30389 38743
rect 30055 38712 30389 38740
rect 30055 38709 30067 38712
rect 30009 38703 30067 38709
rect 30377 38709 30389 38712
rect 30423 38709 30435 38743
rect 30484 38740 30512 38780
rect 30650 38768 30656 38820
rect 30708 38808 30714 38820
rect 30837 38811 30895 38817
rect 30837 38808 30849 38811
rect 30708 38780 30849 38808
rect 30708 38768 30714 38780
rect 30837 38777 30849 38780
rect 30883 38777 30895 38811
rect 30837 38771 30895 38777
rect 31938 38768 31944 38820
rect 31996 38808 32002 38820
rect 32968 38808 32996 38839
rect 33520 38820 33548 38848
rect 33962 38836 33968 38888
rect 34020 38836 34026 38888
rect 34149 38879 34207 38885
rect 34149 38845 34161 38879
rect 34195 38845 34207 38879
rect 34149 38839 34207 38845
rect 31996 38780 32996 38808
rect 31996 38768 32002 38780
rect 33226 38768 33232 38820
rect 33284 38808 33290 38820
rect 33321 38811 33379 38817
rect 33321 38808 33333 38811
rect 33284 38780 33333 38808
rect 33284 38768 33290 38780
rect 33321 38777 33333 38780
rect 33367 38777 33379 38811
rect 33321 38771 33379 38777
rect 33502 38768 33508 38820
rect 33560 38768 33566 38820
rect 33778 38768 33784 38820
rect 33836 38808 33842 38820
rect 34164 38808 34192 38839
rect 33836 38780 34192 38808
rect 33836 38768 33842 38780
rect 34256 38740 34284 38984
rect 35618 38904 35624 38956
rect 35676 38904 35682 38956
rect 35728 38944 35756 38984
rect 36924 38984 37556 39012
rect 36924 38944 36952 38984
rect 37550 38972 37556 38984
rect 37608 38972 37614 39024
rect 37642 38972 37648 39024
rect 37700 38972 37706 39024
rect 37734 38972 37740 39024
rect 37792 39012 37798 39024
rect 37792 38984 38608 39012
rect 37792 38972 37798 38984
rect 35728 38916 36952 38944
rect 37366 38904 37372 38956
rect 37424 38944 37430 38956
rect 38197 38947 38255 38953
rect 38197 38944 38209 38947
rect 37424 38916 38209 38944
rect 37424 38904 37430 38916
rect 38197 38913 38209 38916
rect 38243 38913 38255 38947
rect 38197 38907 38255 38913
rect 35529 38879 35587 38885
rect 35529 38845 35541 38879
rect 35575 38845 35587 38879
rect 35529 38839 35587 38845
rect 30484 38712 34284 38740
rect 30377 38703 30435 38709
rect 34698 38700 34704 38752
rect 34756 38740 34762 38752
rect 34793 38743 34851 38749
rect 34793 38740 34805 38743
rect 34756 38712 34805 38740
rect 34756 38700 34762 38712
rect 34793 38709 34805 38712
rect 34839 38709 34851 38743
rect 34793 38703 34851 38709
rect 34882 38700 34888 38752
rect 34940 38700 34946 38752
rect 35544 38740 35572 38839
rect 37274 38836 37280 38888
rect 37332 38876 37338 38888
rect 38105 38879 38163 38885
rect 38105 38876 38117 38879
rect 37332 38848 38117 38876
rect 37332 38836 37338 38848
rect 38105 38845 38117 38848
rect 38151 38845 38163 38879
rect 38105 38839 38163 38845
rect 38286 38836 38292 38888
rect 38344 38876 38350 38888
rect 38473 38879 38531 38885
rect 38473 38876 38485 38879
rect 38344 38848 38485 38876
rect 38344 38836 38350 38848
rect 38473 38845 38485 38848
rect 38519 38845 38531 38879
rect 38580 38876 38608 38984
rect 39206 38972 39212 39024
rect 39264 39012 39270 39024
rect 39301 39015 39359 39021
rect 39301 39012 39313 39015
rect 39264 38984 39313 39012
rect 39264 38972 39270 38984
rect 39301 38981 39313 38984
rect 39347 38981 39359 39015
rect 39301 38975 39359 38981
rect 39390 38972 39396 39024
rect 39448 39012 39454 39024
rect 40126 39012 40132 39024
rect 39448 38984 40132 39012
rect 39448 38972 39454 38984
rect 40126 38972 40132 38984
rect 40184 38972 40190 39024
rect 40402 38972 40408 39024
rect 40460 39012 40466 39024
rect 40460 38984 40632 39012
rect 40460 38972 40466 38984
rect 39482 38904 39488 38956
rect 39540 38944 39546 38956
rect 39853 38947 39911 38953
rect 39853 38944 39865 38947
rect 39540 38916 39865 38944
rect 39540 38904 39546 38916
rect 39853 38913 39865 38916
rect 39899 38944 39911 38947
rect 40494 38944 40500 38956
rect 39899 38916 40500 38944
rect 39899 38913 39911 38916
rect 39853 38907 39911 38913
rect 40494 38904 40500 38916
rect 40552 38904 40558 38956
rect 40604 38953 40632 38984
rect 47964 38984 50476 39012
rect 40589 38947 40647 38953
rect 40589 38913 40601 38947
rect 40635 38913 40647 38947
rect 40589 38907 40647 38913
rect 40678 38904 40684 38956
rect 40736 38944 40742 38956
rect 40954 38944 40960 38956
rect 40736 38916 40960 38944
rect 40736 38904 40742 38916
rect 40954 38904 40960 38916
rect 41012 38944 41018 38956
rect 41322 38944 41328 38956
rect 41012 38916 41328 38944
rect 41012 38904 41018 38916
rect 41322 38904 41328 38916
rect 41380 38904 41386 38956
rect 41509 38947 41567 38953
rect 41509 38913 41521 38947
rect 41555 38944 41567 38947
rect 42518 38944 42524 38956
rect 41555 38916 42524 38944
rect 41555 38913 41567 38916
rect 41509 38907 41567 38913
rect 39574 38876 39580 38888
rect 38580 38848 39580 38876
rect 38473 38839 38531 38845
rect 39574 38836 39580 38848
rect 39632 38876 39638 38888
rect 39669 38879 39727 38885
rect 39669 38876 39681 38879
rect 39632 38848 39681 38876
rect 39632 38836 39638 38848
rect 39669 38845 39681 38848
rect 39715 38845 39727 38879
rect 39669 38839 39727 38845
rect 39758 38836 39764 38888
rect 39816 38876 39822 38888
rect 41524 38876 41552 38907
rect 42518 38904 42524 38916
rect 42576 38904 42582 38956
rect 43254 38904 43260 38956
rect 43312 38944 43318 38956
rect 43901 38947 43959 38953
rect 43901 38944 43913 38947
rect 43312 38916 43913 38944
rect 43312 38904 43318 38916
rect 43901 38913 43913 38916
rect 43947 38913 43959 38947
rect 43901 38907 43959 38913
rect 44358 38904 44364 38956
rect 44416 38944 44422 38956
rect 45005 38947 45063 38953
rect 45005 38944 45017 38947
rect 44416 38916 45017 38944
rect 44416 38904 44422 38916
rect 45005 38913 45017 38916
rect 45051 38944 45063 38947
rect 47118 38944 47124 38956
rect 45051 38916 47124 38944
rect 45051 38913 45063 38916
rect 45005 38907 45063 38913
rect 47118 38904 47124 38916
rect 47176 38944 47182 38956
rect 47964 38944 47992 38984
rect 47176 38916 47992 38944
rect 47176 38904 47182 38916
rect 48682 38904 48688 38956
rect 48740 38944 48746 38956
rect 49145 38947 49203 38953
rect 49145 38944 49157 38947
rect 48740 38916 49157 38944
rect 48740 38904 48746 38916
rect 49145 38913 49157 38916
rect 49191 38913 49203 38947
rect 49145 38907 49203 38913
rect 49234 38904 49240 38956
rect 49292 38904 49298 38956
rect 50448 38953 50476 38984
rect 50433 38947 50491 38953
rect 50433 38913 50445 38947
rect 50479 38913 50491 38947
rect 50433 38907 50491 38913
rect 53929 38947 53987 38953
rect 53929 38913 53941 38947
rect 53975 38944 53987 38947
rect 55033 38947 55091 38953
rect 55033 38944 55045 38947
rect 53975 38916 55045 38944
rect 53975 38913 53987 38916
rect 53929 38907 53987 38913
rect 55033 38913 55045 38916
rect 55079 38944 55091 38947
rect 56042 38944 56048 38956
rect 55079 38916 56048 38944
rect 55079 38913 55091 38916
rect 55033 38907 55091 38913
rect 56042 38904 56048 38916
rect 56100 38904 56106 38956
rect 56318 38904 56324 38956
rect 56376 38944 56382 38956
rect 57422 38944 57428 38956
rect 56376 38916 57428 38944
rect 56376 38904 56382 38916
rect 57422 38904 57428 38916
rect 57480 38944 57486 38956
rect 58636 38953 58664 39052
rect 60458 39040 60464 39052
rect 60516 39040 60522 39092
rect 58897 39015 58955 39021
rect 58897 38981 58909 39015
rect 58943 39012 58955 39015
rect 59538 39012 59544 39024
rect 58943 38984 59544 39012
rect 58943 38981 58955 38984
rect 58897 38975 58955 38981
rect 59538 38972 59544 38984
rect 59596 38972 59602 39024
rect 58621 38947 58679 38953
rect 58621 38944 58633 38947
rect 57480 38916 58633 38944
rect 57480 38904 57486 38916
rect 58621 38913 58633 38916
rect 58667 38913 58679 38947
rect 58621 38907 58679 38913
rect 59170 38904 59176 38956
rect 59228 38944 59234 38956
rect 59449 38947 59507 38953
rect 59449 38944 59461 38947
rect 59228 38916 59461 38944
rect 59228 38904 59234 38916
rect 59449 38913 59461 38916
rect 59495 38913 59507 38947
rect 59449 38907 59507 38913
rect 59630 38904 59636 38956
rect 59688 38944 59694 38956
rect 60461 38947 60519 38953
rect 60461 38944 60473 38947
rect 59688 38916 60473 38944
rect 59688 38904 59694 38916
rect 60461 38913 60473 38916
rect 60507 38913 60519 38947
rect 60461 38907 60519 38913
rect 39816 38848 41552 38876
rect 39816 38836 39822 38848
rect 43714 38836 43720 38888
rect 43772 38876 43778 38888
rect 45833 38879 45891 38885
rect 45833 38876 45845 38879
rect 43772 38848 45845 38876
rect 43772 38836 43778 38848
rect 45833 38845 45845 38848
rect 45879 38845 45891 38879
rect 45833 38839 45891 38845
rect 46474 38836 46480 38888
rect 46532 38836 46538 38888
rect 47854 38836 47860 38888
rect 47912 38876 47918 38888
rect 48130 38876 48136 38888
rect 47912 38848 48136 38876
rect 47912 38836 47918 38848
rect 48130 38836 48136 38848
rect 48188 38836 48194 38888
rect 48406 38836 48412 38888
rect 48464 38876 48470 38888
rect 49053 38879 49111 38885
rect 49053 38876 49065 38879
rect 48464 38848 49065 38876
rect 48464 38836 48470 38848
rect 49053 38845 49065 38848
rect 49099 38845 49111 38879
rect 49053 38839 49111 38845
rect 51442 38836 51448 38888
rect 51500 38836 51506 38888
rect 57790 38836 57796 38888
rect 57848 38876 57854 38888
rect 58529 38879 58587 38885
rect 58529 38876 58541 38879
rect 57848 38848 58541 38876
rect 57848 38836 57854 38848
rect 58529 38845 58541 38848
rect 58575 38845 58587 38879
rect 58529 38839 58587 38845
rect 59265 38879 59323 38885
rect 59265 38845 59277 38879
rect 59311 38876 59323 38879
rect 60274 38876 60280 38888
rect 59311 38848 60280 38876
rect 59311 38845 59323 38848
rect 59265 38839 59323 38845
rect 60274 38836 60280 38848
rect 60332 38836 60338 38888
rect 35894 38768 35900 38820
rect 35952 38768 35958 38820
rect 37182 38808 37188 38820
rect 37122 38780 37188 38808
rect 37182 38768 37188 38780
rect 37240 38768 37246 38820
rect 37458 38768 37464 38820
rect 37516 38808 37522 38820
rect 38013 38811 38071 38817
rect 38013 38808 38025 38811
rect 37516 38780 38025 38808
rect 37516 38768 37522 38780
rect 38013 38777 38025 38780
rect 38059 38777 38071 38811
rect 38013 38771 38071 38777
rect 38120 38780 39804 38808
rect 36814 38740 36820 38752
rect 35544 38712 36820 38740
rect 36814 38700 36820 38712
rect 36872 38700 36878 38752
rect 37366 38700 37372 38752
rect 37424 38740 37430 38752
rect 38120 38740 38148 38780
rect 37424 38712 38148 38740
rect 37424 38700 37430 38712
rect 39114 38700 39120 38752
rect 39172 38700 39178 38752
rect 39776 38749 39804 38780
rect 41782 38768 41788 38820
rect 41840 38768 41846 38820
rect 44821 38811 44879 38817
rect 41892 38780 42274 38808
rect 39761 38743 39819 38749
rect 39761 38709 39773 38743
rect 39807 38709 39819 38743
rect 39761 38703 39819 38709
rect 40126 38700 40132 38752
rect 40184 38700 40190 38752
rect 40494 38700 40500 38752
rect 40552 38700 40558 38752
rect 41046 38700 41052 38752
rect 41104 38740 41110 38752
rect 41892 38740 41920 38780
rect 44821 38777 44833 38811
rect 44867 38808 44879 38811
rect 45646 38808 45652 38820
rect 44867 38780 45652 38808
rect 44867 38777 44879 38780
rect 44821 38771 44879 38777
rect 45646 38768 45652 38780
rect 45704 38768 45710 38820
rect 47578 38768 47584 38820
rect 47636 38768 47642 38820
rect 50249 38811 50307 38817
rect 50249 38777 50261 38811
rect 50295 38808 50307 38811
rect 50893 38811 50951 38817
rect 50893 38808 50905 38811
rect 50295 38780 50905 38808
rect 50295 38777 50307 38780
rect 50249 38771 50307 38777
rect 50893 38777 50905 38780
rect 50939 38777 50951 38811
rect 50893 38771 50951 38777
rect 53006 38768 53012 38820
rect 53064 38768 53070 38820
rect 53650 38768 53656 38820
rect 53708 38768 53714 38820
rect 55306 38768 55312 38820
rect 55364 38768 55370 38820
rect 55766 38808 55772 38820
rect 55600 38780 55772 38808
rect 41104 38712 41920 38740
rect 41104 38700 41110 38712
rect 44082 38700 44088 38752
rect 44140 38740 44146 38752
rect 44453 38743 44511 38749
rect 44453 38740 44465 38743
rect 44140 38712 44465 38740
rect 44140 38700 44146 38712
rect 44453 38709 44465 38712
rect 44499 38709 44511 38743
rect 44453 38703 44511 38709
rect 44910 38700 44916 38752
rect 44968 38700 44974 38752
rect 46934 38700 46940 38752
rect 46992 38740 46998 38752
rect 47854 38740 47860 38752
rect 46992 38712 47860 38740
rect 46992 38700 46998 38712
rect 47854 38700 47860 38712
rect 47912 38700 47918 38752
rect 49878 38700 49884 38752
rect 49936 38700 49942 38752
rect 50338 38700 50344 38752
rect 50396 38700 50402 38752
rect 52181 38743 52239 38749
rect 52181 38709 52193 38743
rect 52227 38740 52239 38743
rect 53558 38740 53564 38752
rect 52227 38712 53564 38740
rect 52227 38709 52239 38712
rect 52181 38703 52239 38709
rect 53558 38700 53564 38712
rect 53616 38700 53622 38752
rect 55214 38700 55220 38752
rect 55272 38740 55278 38752
rect 55600 38740 55628 38780
rect 55766 38768 55772 38780
rect 55824 38768 55830 38820
rect 58437 38811 58495 38817
rect 58437 38777 58449 38811
rect 58483 38808 58495 38811
rect 59909 38811 59967 38817
rect 59909 38808 59921 38811
rect 58483 38780 59921 38808
rect 58483 38777 58495 38780
rect 58437 38771 58495 38777
rect 59909 38777 59921 38780
rect 59955 38777 59967 38811
rect 59909 38771 59967 38777
rect 55272 38712 55628 38740
rect 55272 38700 55278 38712
rect 56778 38700 56784 38752
rect 56836 38700 56842 38752
rect 58069 38743 58127 38749
rect 58069 38709 58081 38743
rect 58115 38740 58127 38743
rect 58158 38740 58164 38752
rect 58115 38712 58164 38740
rect 58115 38709 58127 38712
rect 58069 38703 58127 38709
rect 58158 38700 58164 38712
rect 58216 38700 58222 38752
rect 59170 38700 59176 38752
rect 59228 38740 59234 38752
rect 59357 38743 59415 38749
rect 59357 38740 59369 38743
rect 59228 38712 59369 38740
rect 59228 38700 59234 38712
rect 59357 38709 59369 38712
rect 59403 38709 59415 38743
rect 59357 38703 59415 38709
rect 552 38650 66424 38672
rect 552 38598 2918 38650
rect 2970 38598 2982 38650
rect 3034 38598 3046 38650
rect 3098 38598 3110 38650
rect 3162 38598 3174 38650
rect 3226 38598 50918 38650
rect 50970 38598 50982 38650
rect 51034 38598 51046 38650
rect 51098 38598 51110 38650
rect 51162 38598 51174 38650
rect 51226 38598 66424 38650
rect 552 38576 66424 38598
rect 8386 38536 8392 38548
rect 7116 38508 8392 38536
rect 7116 38409 7144 38508
rect 8386 38496 8392 38508
rect 8444 38496 8450 38548
rect 8662 38496 8668 38548
rect 8720 38536 8726 38548
rect 8846 38536 8852 38548
rect 8720 38508 8852 38536
rect 8720 38496 8726 38508
rect 8846 38496 8852 38508
rect 8904 38496 8910 38548
rect 9122 38496 9128 38548
rect 9180 38536 9186 38548
rect 9217 38539 9275 38545
rect 9217 38536 9229 38539
rect 9180 38508 9229 38536
rect 9180 38496 9186 38508
rect 9217 38505 9229 38508
rect 9263 38505 9275 38539
rect 9217 38499 9275 38505
rect 9490 38496 9496 38548
rect 9548 38536 9554 38548
rect 9585 38539 9643 38545
rect 9585 38536 9597 38539
rect 9548 38508 9597 38536
rect 9548 38496 9554 38508
rect 9585 38505 9597 38508
rect 9631 38505 9643 38539
rect 9585 38499 9643 38505
rect 10781 38539 10839 38545
rect 10781 38505 10793 38539
rect 10827 38536 10839 38539
rect 10870 38536 10876 38548
rect 10827 38508 10876 38536
rect 10827 38505 10839 38508
rect 10781 38499 10839 38505
rect 10870 38496 10876 38508
rect 10928 38496 10934 38548
rect 11238 38496 11244 38548
rect 11296 38536 11302 38548
rect 11296 38508 13584 38536
rect 11296 38496 11302 38508
rect 10413 38471 10471 38477
rect 10413 38437 10425 38471
rect 10459 38468 10471 38471
rect 11977 38471 12035 38477
rect 11977 38468 11989 38471
rect 10459 38440 11989 38468
rect 10459 38437 10471 38440
rect 10413 38431 10471 38437
rect 11977 38437 11989 38440
rect 12023 38437 12035 38471
rect 11977 38431 12035 38437
rect 7101 38403 7159 38409
rect 7101 38369 7113 38403
rect 7147 38369 7159 38403
rect 9950 38400 9956 38412
rect 8510 38372 9956 38400
rect 7101 38363 7159 38369
rect 9950 38360 9956 38372
rect 10008 38360 10014 38412
rect 11238 38400 11244 38412
rect 10152 38372 11244 38400
rect 7377 38335 7435 38341
rect 7377 38301 7389 38335
rect 7423 38332 7435 38335
rect 7466 38332 7472 38344
rect 7423 38304 7472 38332
rect 7423 38301 7435 38304
rect 7377 38295 7435 38301
rect 7466 38292 7472 38304
rect 7524 38292 7530 38344
rect 9674 38292 9680 38344
rect 9732 38292 9738 38344
rect 9861 38335 9919 38341
rect 9861 38301 9873 38335
rect 9907 38332 9919 38335
rect 10152 38332 10180 38372
rect 11238 38360 11244 38372
rect 11296 38360 11302 38412
rect 11517 38403 11575 38409
rect 11517 38369 11529 38403
rect 11563 38400 11575 38403
rect 12342 38400 12348 38412
rect 11563 38372 12348 38400
rect 11563 38369 11575 38372
rect 11517 38363 11575 38369
rect 12342 38360 12348 38372
rect 12400 38400 12406 38412
rect 12529 38403 12587 38409
rect 12529 38400 12541 38403
rect 12400 38372 12541 38400
rect 12400 38360 12406 38372
rect 12529 38369 12541 38372
rect 12575 38369 12587 38403
rect 13556 38400 13584 38508
rect 13630 38496 13636 38548
rect 13688 38536 13694 38548
rect 14001 38539 14059 38545
rect 14001 38536 14013 38539
rect 13688 38508 14013 38536
rect 13688 38496 13694 38508
rect 14001 38505 14013 38508
rect 14047 38505 14059 38539
rect 14001 38499 14059 38505
rect 14458 38496 14464 38548
rect 14516 38496 14522 38548
rect 15657 38539 15715 38545
rect 15657 38505 15669 38539
rect 15703 38536 15715 38539
rect 16482 38536 16488 38548
rect 15703 38508 16488 38536
rect 15703 38505 15715 38508
rect 15657 38499 15715 38505
rect 16482 38496 16488 38508
rect 16540 38496 16546 38548
rect 19334 38496 19340 38548
rect 19392 38536 19398 38548
rect 20165 38539 20223 38545
rect 20165 38536 20177 38539
rect 19392 38508 20177 38536
rect 19392 38496 19398 38508
rect 20165 38505 20177 38508
rect 20211 38505 20223 38539
rect 20165 38499 20223 38505
rect 20530 38496 20536 38548
rect 20588 38496 20594 38548
rect 21634 38496 21640 38548
rect 21692 38496 21698 38548
rect 22094 38536 22100 38548
rect 21744 38508 22100 38536
rect 14093 38471 14151 38477
rect 14093 38437 14105 38471
rect 14139 38468 14151 38471
rect 15194 38468 15200 38480
rect 14139 38440 15200 38468
rect 14139 38437 14151 38440
rect 14093 38431 14151 38437
rect 15194 38428 15200 38440
rect 15252 38428 15258 38480
rect 15470 38428 15476 38480
rect 15528 38468 15534 38480
rect 15528 38440 17632 38468
rect 15528 38428 15534 38440
rect 17604 38412 17632 38440
rect 19242 38428 19248 38480
rect 19300 38468 19306 38480
rect 21744 38468 21772 38508
rect 22094 38496 22100 38508
rect 22152 38496 22158 38548
rect 22186 38496 22192 38548
rect 22244 38536 22250 38548
rect 23109 38539 23167 38545
rect 23109 38536 23121 38539
rect 22244 38508 23121 38536
rect 22244 38496 22250 38508
rect 23109 38505 23121 38508
rect 23155 38505 23167 38539
rect 23109 38499 23167 38505
rect 23477 38539 23535 38545
rect 23477 38505 23489 38539
rect 23523 38536 23535 38539
rect 23842 38536 23848 38548
rect 23523 38508 23848 38536
rect 23523 38505 23535 38508
rect 23477 38499 23535 38505
rect 23842 38496 23848 38508
rect 23900 38496 23906 38548
rect 24578 38496 24584 38548
rect 24636 38536 24642 38548
rect 24636 38508 25728 38536
rect 24636 38496 24642 38508
rect 19300 38440 21772 38468
rect 19300 38428 19306 38440
rect 21910 38428 21916 38480
rect 21968 38468 21974 38480
rect 21968 38440 24164 38468
rect 21968 38428 21974 38440
rect 13556 38372 13952 38400
rect 12529 38363 12587 38369
rect 9907 38304 10180 38332
rect 10229 38335 10287 38341
rect 9907 38301 9919 38304
rect 9861 38295 9919 38301
rect 10229 38301 10241 38335
rect 10275 38301 10287 38335
rect 10229 38295 10287 38301
rect 10321 38335 10379 38341
rect 10321 38301 10333 38335
rect 10367 38332 10379 38335
rect 11330 38332 11336 38344
rect 10367 38304 11336 38332
rect 10367 38301 10379 38304
rect 10321 38295 10379 38301
rect 9306 38224 9312 38276
rect 9364 38264 9370 38276
rect 10244 38264 10272 38295
rect 11330 38292 11336 38304
rect 11388 38292 11394 38344
rect 11609 38335 11667 38341
rect 11609 38301 11621 38335
rect 11655 38301 11667 38335
rect 11609 38295 11667 38301
rect 11793 38335 11851 38341
rect 11793 38301 11805 38335
rect 11839 38332 11851 38335
rect 12802 38332 12808 38344
rect 11839 38304 12808 38332
rect 11839 38301 11851 38304
rect 11793 38295 11851 38301
rect 11624 38264 11652 38295
rect 12802 38292 12808 38304
rect 12860 38332 12866 38344
rect 13722 38332 13728 38344
rect 12860 38304 13728 38332
rect 12860 38292 12866 38304
rect 13722 38292 13728 38304
rect 13780 38292 13786 38344
rect 13924 38341 13952 38372
rect 15286 38360 15292 38412
rect 15344 38400 15350 38412
rect 15565 38403 15623 38409
rect 15565 38400 15577 38403
rect 15344 38372 15577 38400
rect 15344 38360 15350 38372
rect 15565 38369 15577 38372
rect 15611 38369 15623 38403
rect 15565 38363 15623 38369
rect 15672 38372 16344 38400
rect 13909 38335 13967 38341
rect 13909 38301 13921 38335
rect 13955 38332 13967 38335
rect 15672 38332 15700 38372
rect 13955 38304 15700 38332
rect 15841 38335 15899 38341
rect 13955 38301 13967 38304
rect 13909 38295 13967 38301
rect 15841 38301 15853 38335
rect 15887 38332 15899 38335
rect 15887 38304 16068 38332
rect 15887 38301 15899 38304
rect 15841 38295 15899 38301
rect 12618 38264 12624 38276
rect 9364 38236 11284 38264
rect 11624 38236 12624 38264
rect 9364 38224 9370 38236
rect 10962 38156 10968 38208
rect 11020 38196 11026 38208
rect 11149 38199 11207 38205
rect 11149 38196 11161 38199
rect 11020 38168 11161 38196
rect 11020 38156 11026 38168
rect 11149 38165 11161 38168
rect 11195 38165 11207 38199
rect 11256 38196 11284 38236
rect 12618 38224 12624 38236
rect 12676 38224 12682 38276
rect 14550 38224 14556 38276
rect 14608 38264 14614 38276
rect 16040 38264 16068 38304
rect 16316 38264 16344 38372
rect 16482 38360 16488 38412
rect 16540 38360 16546 38412
rect 17586 38360 17592 38412
rect 17644 38360 17650 38412
rect 17678 38360 17684 38412
rect 17736 38400 17742 38412
rect 17736 38372 22416 38400
rect 17736 38360 17742 38372
rect 16390 38292 16396 38344
rect 16448 38332 16454 38344
rect 16577 38335 16635 38341
rect 16577 38332 16589 38335
rect 16448 38304 16589 38332
rect 16448 38292 16454 38304
rect 16577 38301 16589 38304
rect 16623 38301 16635 38335
rect 16577 38295 16635 38301
rect 16669 38335 16727 38341
rect 16669 38301 16681 38335
rect 16715 38301 16727 38335
rect 16669 38295 16727 38301
rect 16684 38264 16712 38295
rect 18782 38292 18788 38344
rect 18840 38332 18846 38344
rect 19889 38335 19947 38341
rect 19889 38332 19901 38335
rect 18840 38304 19901 38332
rect 18840 38292 18846 38304
rect 19889 38301 19901 38304
rect 19935 38301 19947 38335
rect 19889 38295 19947 38301
rect 20073 38335 20131 38341
rect 20073 38301 20085 38335
rect 20119 38301 20131 38335
rect 20073 38295 20131 38301
rect 20180 38304 21588 38332
rect 14608 38236 15332 38264
rect 16040 38236 16252 38264
rect 16316 38236 16712 38264
rect 14608 38224 14614 38236
rect 14366 38196 14372 38208
rect 11256 38168 14372 38196
rect 11149 38159 11207 38165
rect 14366 38156 14372 38168
rect 14424 38156 14430 38208
rect 15194 38156 15200 38208
rect 15252 38156 15258 38208
rect 15304 38196 15332 38236
rect 16117 38199 16175 38205
rect 16117 38196 16129 38199
rect 15304 38168 16129 38196
rect 16117 38165 16129 38168
rect 16163 38165 16175 38199
rect 16224 38196 16252 38236
rect 17862 38224 17868 38276
rect 17920 38264 17926 38276
rect 20088 38264 20116 38295
rect 17920 38236 20116 38264
rect 17920 38224 17926 38236
rect 19242 38196 19248 38208
rect 16224 38168 19248 38196
rect 16117 38159 16175 38165
rect 19242 38156 19248 38168
rect 19300 38156 19306 38208
rect 19334 38156 19340 38208
rect 19392 38196 19398 38208
rect 20180 38196 20208 38304
rect 20714 38224 20720 38276
rect 20772 38264 20778 38276
rect 21450 38264 21456 38276
rect 20772 38236 21456 38264
rect 20772 38224 20778 38236
rect 21450 38224 21456 38236
rect 21508 38224 21514 38276
rect 21560 38264 21588 38304
rect 21726 38292 21732 38344
rect 21784 38292 21790 38344
rect 21913 38335 21971 38341
rect 21913 38301 21925 38335
rect 21959 38301 21971 38335
rect 21913 38295 21971 38301
rect 21928 38264 21956 38295
rect 22189 38267 22247 38273
rect 22189 38264 22201 38267
rect 21560 38236 22201 38264
rect 22189 38233 22201 38236
rect 22235 38233 22247 38267
rect 22189 38227 22247 38233
rect 19392 38168 20208 38196
rect 19392 38156 19398 38168
rect 20898 38156 20904 38208
rect 20956 38196 20962 38208
rect 21269 38199 21327 38205
rect 21269 38196 21281 38199
rect 20956 38168 21281 38196
rect 20956 38156 20962 38168
rect 21269 38165 21281 38168
rect 21315 38165 21327 38199
rect 22388 38196 22416 38372
rect 22462 38360 22468 38412
rect 22520 38360 22526 38412
rect 24136 38409 24164 38440
rect 25038 38428 25044 38480
rect 25096 38428 25102 38480
rect 25700 38468 25728 38508
rect 26234 38496 26240 38548
rect 26292 38536 26298 38548
rect 29546 38536 29552 38548
rect 26292 38508 29552 38536
rect 26292 38496 26298 38508
rect 26970 38468 26976 38480
rect 25700 38440 26976 38468
rect 26970 38428 26976 38440
rect 27028 38428 27034 38480
rect 27341 38471 27399 38477
rect 27341 38437 27353 38471
rect 27387 38468 27399 38471
rect 27614 38468 27620 38480
rect 27387 38440 27620 38468
rect 27387 38437 27399 38440
rect 27341 38431 27399 38437
rect 27614 38428 27620 38440
rect 27672 38428 27678 38480
rect 24121 38403 24179 38409
rect 24121 38369 24133 38403
rect 24167 38369 24179 38403
rect 24121 38363 24179 38369
rect 28442 38360 28448 38412
rect 28500 38360 28506 38412
rect 28920 38409 28948 38508
rect 29546 38496 29552 38508
rect 29604 38496 29610 38548
rect 29914 38496 29920 38548
rect 29972 38536 29978 38548
rect 30745 38539 30803 38545
rect 30745 38536 30757 38539
rect 29972 38508 30757 38536
rect 29972 38496 29978 38508
rect 30745 38505 30757 38508
rect 30791 38505 30803 38539
rect 30745 38499 30803 38505
rect 33134 38496 33140 38548
rect 33192 38536 33198 38548
rect 33192 38508 34836 38536
rect 33192 38496 33198 38508
rect 29178 38428 29184 38480
rect 29236 38428 29242 38480
rect 31202 38468 31208 38480
rect 30406 38440 31208 38468
rect 31202 38428 31208 38440
rect 31260 38468 31266 38480
rect 31386 38468 31392 38480
rect 31260 38440 31392 38468
rect 31260 38428 31266 38440
rect 31386 38428 31392 38440
rect 31444 38428 31450 38480
rect 33870 38428 33876 38480
rect 33928 38428 33934 38480
rect 34808 38468 34836 38508
rect 34882 38496 34888 38548
rect 34940 38536 34946 38548
rect 35345 38539 35403 38545
rect 35345 38536 35357 38539
rect 34940 38508 35357 38536
rect 34940 38496 34946 38508
rect 35345 38505 35357 38508
rect 35391 38505 35403 38539
rect 35345 38499 35403 38505
rect 35437 38539 35495 38545
rect 35437 38505 35449 38539
rect 35483 38536 35495 38539
rect 35805 38539 35863 38545
rect 35805 38536 35817 38539
rect 35483 38508 35817 38536
rect 35483 38505 35495 38508
rect 35437 38499 35495 38505
rect 35805 38505 35817 38508
rect 35851 38505 35863 38539
rect 35805 38499 35863 38505
rect 35894 38496 35900 38548
rect 35952 38536 35958 38548
rect 36725 38539 36783 38545
rect 36725 38536 36737 38539
rect 35952 38508 36737 38536
rect 35952 38496 35958 38508
rect 36725 38505 36737 38508
rect 36771 38505 36783 38539
rect 36725 38499 36783 38505
rect 36814 38496 36820 38548
rect 36872 38536 36878 38548
rect 37093 38539 37151 38545
rect 37093 38536 37105 38539
rect 36872 38508 37105 38536
rect 36872 38496 36878 38508
rect 37093 38505 37105 38508
rect 37139 38505 37151 38539
rect 37093 38499 37151 38505
rect 38197 38539 38255 38545
rect 38197 38505 38209 38539
rect 38243 38536 38255 38539
rect 38286 38536 38292 38548
rect 38243 38508 38292 38536
rect 38243 38505 38255 38508
rect 38197 38499 38255 38505
rect 38286 38496 38292 38508
rect 38344 38496 38350 38548
rect 38396 38508 39988 38536
rect 34808 38440 35020 38468
rect 28905 38403 28963 38409
rect 28905 38369 28917 38403
rect 28951 38369 28963 38403
rect 28905 38363 28963 38369
rect 30576 38372 31432 38400
rect 23566 38292 23572 38344
rect 23624 38292 23630 38344
rect 23753 38335 23811 38341
rect 23753 38301 23765 38335
rect 23799 38332 23811 38335
rect 24026 38332 24032 38344
rect 23799 38304 24032 38332
rect 23799 38301 23811 38304
rect 23753 38295 23811 38301
rect 24026 38292 24032 38304
rect 24084 38292 24090 38344
rect 24397 38335 24455 38341
rect 24397 38301 24409 38335
rect 24443 38332 24455 38335
rect 25682 38332 25688 38344
rect 24443 38304 25688 38332
rect 24443 38301 24455 38304
rect 24397 38295 24455 38301
rect 25682 38292 25688 38304
rect 25740 38292 25746 38344
rect 27062 38292 27068 38344
rect 27120 38292 27126 38344
rect 30576 38332 30604 38372
rect 27172 38304 30604 38332
rect 30653 38335 30711 38341
rect 27172 38264 27200 38304
rect 30653 38301 30665 38335
rect 30699 38332 30711 38335
rect 30742 38332 30748 38344
rect 30699 38304 30748 38332
rect 30699 38301 30711 38304
rect 30653 38295 30711 38301
rect 30742 38292 30748 38304
rect 30800 38332 30806 38344
rect 31297 38335 31355 38341
rect 31297 38332 31309 38335
rect 30800 38304 31309 38332
rect 30800 38292 30806 38304
rect 31297 38301 31309 38304
rect 31343 38301 31355 38335
rect 31404 38332 31432 38372
rect 32950 38360 32956 38412
rect 33008 38400 33014 38412
rect 33226 38400 33232 38412
rect 33008 38372 33232 38400
rect 33008 38360 33014 38372
rect 33226 38360 33232 38372
rect 33284 38360 33290 38412
rect 34882 38360 34888 38412
rect 34940 38360 34946 38412
rect 34992 38400 35020 38440
rect 36262 38428 36268 38480
rect 36320 38428 36326 38480
rect 36173 38403 36231 38409
rect 36173 38400 36185 38403
rect 34992 38372 36185 38400
rect 36173 38369 36185 38372
rect 36219 38400 36231 38403
rect 37185 38403 37243 38409
rect 37185 38400 37197 38403
rect 36219 38372 37197 38400
rect 36219 38369 36231 38372
rect 36173 38363 36231 38369
rect 37185 38369 37197 38372
rect 37231 38400 37243 38403
rect 37366 38400 37372 38412
rect 37231 38372 37372 38400
rect 37231 38369 37243 38372
rect 37185 38363 37243 38369
rect 37366 38360 37372 38372
rect 37424 38360 37430 38412
rect 34609 38335 34667 38341
rect 31404 38304 33640 38332
rect 31297 38295 31355 38301
rect 25424 38236 27200 38264
rect 25424 38196 25452 38236
rect 28350 38224 28356 38276
rect 28408 38264 28414 38276
rect 28408 38236 28948 38264
rect 28408 38224 28414 38236
rect 22388 38168 25452 38196
rect 21269 38159 21327 38165
rect 25866 38156 25872 38208
rect 25924 38196 25930 38208
rect 27522 38196 27528 38208
rect 25924 38168 27528 38196
rect 25924 38156 25930 38168
rect 27522 38156 27528 38168
rect 27580 38156 27586 38208
rect 28810 38156 28816 38208
rect 28868 38156 28874 38208
rect 28920 38196 28948 38236
rect 32950 38196 32956 38208
rect 28920 38168 32956 38196
rect 32950 38156 32956 38168
rect 33008 38156 33014 38208
rect 33137 38199 33195 38205
rect 33137 38165 33149 38199
rect 33183 38196 33195 38199
rect 33226 38196 33232 38208
rect 33183 38168 33232 38196
rect 33183 38165 33195 38168
rect 33137 38159 33195 38165
rect 33226 38156 33232 38168
rect 33284 38156 33290 38208
rect 33612 38196 33640 38304
rect 34609 38301 34621 38335
rect 34655 38332 34667 38335
rect 35158 38332 35164 38344
rect 34655 38304 34836 38332
rect 34655 38301 34667 38304
rect 34609 38295 34667 38301
rect 34808 38264 34836 38304
rect 35084 38304 35164 38332
rect 34882 38264 34888 38276
rect 34808 38236 34888 38264
rect 34882 38224 34888 38236
rect 34940 38224 34946 38276
rect 34977 38267 35035 38273
rect 34977 38233 34989 38267
rect 35023 38264 35035 38267
rect 35084 38264 35112 38304
rect 35158 38292 35164 38304
rect 35216 38292 35222 38344
rect 35434 38292 35440 38344
rect 35492 38332 35498 38344
rect 35529 38335 35587 38341
rect 35529 38332 35541 38335
rect 35492 38304 35541 38332
rect 35492 38292 35498 38304
rect 35529 38301 35541 38304
rect 35575 38301 35587 38335
rect 35529 38295 35587 38301
rect 35710 38292 35716 38344
rect 35768 38332 35774 38344
rect 36357 38335 36415 38341
rect 36357 38332 36369 38335
rect 35768 38304 36369 38332
rect 35768 38292 35774 38304
rect 36357 38301 36369 38304
rect 36403 38301 36415 38335
rect 36357 38295 36415 38301
rect 37277 38335 37335 38341
rect 37277 38301 37289 38335
rect 37323 38332 37335 38335
rect 38396 38332 38424 38508
rect 39206 38428 39212 38480
rect 39264 38468 39270 38480
rect 39666 38468 39672 38480
rect 39264 38440 39672 38468
rect 39264 38428 39270 38440
rect 39666 38428 39672 38440
rect 39724 38428 39730 38480
rect 39960 38468 39988 38508
rect 40034 38496 40040 38548
rect 40092 38536 40098 38548
rect 40405 38539 40463 38545
rect 40405 38536 40417 38539
rect 40092 38508 40417 38536
rect 40092 38496 40098 38508
rect 40405 38505 40417 38508
rect 40451 38505 40463 38539
rect 40405 38499 40463 38505
rect 40865 38539 40923 38545
rect 40865 38505 40877 38539
rect 40911 38536 40923 38539
rect 41230 38536 41236 38548
rect 40911 38508 41236 38536
rect 40911 38505 40923 38508
rect 40865 38499 40923 38505
rect 41230 38496 41236 38508
rect 41288 38496 41294 38548
rect 42518 38496 42524 38548
rect 42576 38536 42582 38548
rect 44818 38536 44824 38548
rect 42576 38508 44824 38536
rect 42576 38496 42582 38508
rect 40218 38468 40224 38480
rect 39960 38440 40224 38468
rect 40218 38428 40224 38440
rect 40276 38468 40282 38480
rect 41138 38468 41144 38480
rect 40276 38440 41144 38468
rect 40276 38428 40282 38440
rect 41138 38428 41144 38440
rect 41196 38428 41202 38480
rect 43438 38428 43444 38480
rect 43496 38428 43502 38480
rect 40773 38403 40831 38409
rect 40773 38369 40785 38403
rect 40819 38400 40831 38403
rect 41230 38400 41236 38412
rect 40819 38372 41236 38400
rect 40819 38369 40831 38372
rect 40773 38363 40831 38369
rect 41230 38360 41236 38372
rect 41288 38360 41294 38412
rect 41322 38360 41328 38412
rect 41380 38400 41386 38412
rect 43824 38409 43852 38508
rect 44818 38496 44824 38508
rect 44876 38496 44882 38548
rect 45646 38496 45652 38548
rect 45704 38496 45710 38548
rect 47394 38496 47400 38548
rect 47452 38496 47458 38548
rect 47578 38496 47584 38548
rect 47636 38536 47642 38548
rect 47765 38539 47823 38545
rect 47765 38536 47777 38539
rect 47636 38508 47777 38536
rect 47636 38496 47642 38508
rect 47765 38505 47777 38508
rect 47811 38505 47823 38539
rect 47765 38499 47823 38505
rect 48409 38539 48467 38545
rect 48409 38505 48421 38539
rect 48455 38536 48467 38539
rect 48682 38536 48688 38548
rect 48455 38508 48688 38536
rect 48455 38505 48467 38508
rect 48409 38499 48467 38505
rect 48682 38496 48688 38508
rect 48740 38496 48746 38548
rect 48774 38496 48780 38548
rect 48832 38496 48838 38548
rect 48869 38539 48927 38545
rect 48869 38505 48881 38539
rect 48915 38536 48927 38539
rect 51442 38536 51448 38548
rect 48915 38508 51448 38536
rect 48915 38505 48927 38508
rect 48869 38499 48927 38505
rect 51442 38496 51448 38508
rect 51500 38496 51506 38548
rect 53190 38496 53196 38548
rect 53248 38536 53254 38548
rect 53285 38539 53343 38545
rect 53285 38536 53297 38539
rect 53248 38508 53297 38536
rect 53248 38496 53254 38508
rect 53285 38505 53297 38508
rect 53331 38505 53343 38539
rect 53285 38499 53343 38505
rect 53650 38496 53656 38548
rect 53708 38496 53714 38548
rect 59998 38536 60004 38548
rect 53944 38508 60004 38536
rect 44082 38428 44088 38480
rect 44140 38428 44146 38480
rect 47854 38428 47860 38480
rect 47912 38468 47918 38480
rect 47912 38440 49648 38468
rect 47912 38428 47918 38440
rect 49620 38409 49648 38440
rect 49878 38428 49884 38480
rect 49936 38428 49942 38480
rect 49970 38428 49976 38480
rect 50028 38468 50034 38480
rect 50028 38440 50370 38468
rect 50028 38428 50034 38440
rect 51166 38428 51172 38480
rect 51224 38468 51230 38480
rect 53944 38468 53972 38508
rect 59998 38496 60004 38508
rect 60056 38496 60062 38548
rect 60277 38539 60335 38545
rect 60277 38505 60289 38539
rect 60323 38536 60335 38539
rect 60366 38536 60372 38548
rect 60323 38508 60372 38536
rect 60323 38505 60335 38508
rect 60277 38499 60335 38505
rect 60366 38496 60372 38508
rect 60424 38496 60430 38548
rect 51224 38440 53144 38468
rect 51224 38428 51230 38440
rect 43809 38403 43867 38409
rect 41380 38372 42366 38400
rect 41380 38360 41386 38372
rect 43809 38369 43821 38403
rect 43855 38369 43867 38403
rect 49605 38403 49663 38409
rect 45218 38372 45324 38400
rect 43809 38363 43867 38369
rect 45296 38344 45324 38372
rect 49605 38369 49617 38403
rect 49651 38369 49663 38403
rect 49605 38363 49663 38369
rect 51184 38372 52868 38400
rect 39206 38332 39212 38344
rect 37323 38304 38424 38332
rect 38488 38304 39212 38332
rect 37323 38301 37335 38304
rect 37277 38295 37335 38301
rect 35023 38236 35112 38264
rect 35023 38233 35035 38236
rect 34977 38227 35035 38233
rect 37182 38224 37188 38276
rect 37240 38264 37246 38276
rect 38488 38264 38516 38304
rect 39206 38292 39212 38304
rect 39264 38292 39270 38344
rect 39298 38292 39304 38344
rect 39356 38332 39362 38344
rect 39669 38335 39727 38341
rect 39669 38332 39681 38335
rect 39356 38304 39681 38332
rect 39356 38292 39362 38304
rect 39669 38301 39681 38304
rect 39715 38301 39727 38335
rect 39669 38295 39727 38301
rect 39942 38292 39948 38344
rect 40000 38292 40006 38344
rect 41049 38335 41107 38341
rect 41049 38301 41061 38335
rect 41095 38332 41107 38335
rect 41874 38332 41880 38344
rect 41095 38304 41880 38332
rect 41095 38301 41107 38304
rect 41049 38295 41107 38301
rect 41874 38292 41880 38304
rect 41932 38292 41938 38344
rect 43714 38292 43720 38344
rect 43772 38292 43778 38344
rect 45278 38292 45284 38344
rect 45336 38292 45342 38344
rect 45557 38335 45615 38341
rect 45557 38301 45569 38335
rect 45603 38332 45615 38335
rect 45646 38332 45652 38344
rect 45603 38304 45652 38332
rect 45603 38301 45615 38304
rect 45557 38295 45615 38301
rect 45646 38292 45652 38304
rect 45704 38332 45710 38344
rect 46201 38335 46259 38341
rect 46201 38332 46213 38335
rect 45704 38304 46213 38332
rect 45704 38292 45710 38304
rect 46201 38301 46213 38304
rect 46247 38301 46259 38335
rect 46201 38295 46259 38301
rect 47118 38292 47124 38344
rect 47176 38292 47182 38344
rect 47305 38335 47363 38341
rect 47305 38301 47317 38335
rect 47351 38332 47363 38335
rect 47762 38332 47768 38344
rect 47351 38304 47768 38332
rect 47351 38301 47363 38304
rect 47305 38295 47363 38301
rect 47762 38292 47768 38304
rect 47820 38292 47826 38344
rect 48590 38292 48596 38344
rect 48648 38332 48654 38344
rect 48961 38335 49019 38341
rect 48961 38332 48973 38335
rect 48648 38304 48973 38332
rect 48648 38292 48654 38304
rect 48961 38301 48973 38304
rect 49007 38301 49019 38335
rect 51074 38332 51080 38344
rect 48961 38295 49019 38301
rect 49712 38304 51080 38332
rect 37240 38236 38516 38264
rect 37240 38224 37246 38236
rect 41690 38224 41696 38276
rect 41748 38264 41754 38276
rect 41748 38236 42472 38264
rect 41748 38224 41754 38236
rect 41046 38196 41052 38208
rect 33612 38168 41052 38196
rect 41046 38156 41052 38168
rect 41104 38156 41110 38208
rect 41966 38156 41972 38208
rect 42024 38156 42030 38208
rect 42444 38196 42472 38236
rect 45094 38224 45100 38276
rect 45152 38264 45158 38276
rect 49712 38264 49740 38304
rect 51074 38292 51080 38304
rect 51132 38292 51138 38344
rect 45152 38236 49740 38264
rect 45152 38224 45158 38236
rect 43714 38196 43720 38208
rect 42444 38168 43720 38196
rect 43714 38156 43720 38168
rect 43772 38156 43778 38208
rect 44726 38156 44732 38208
rect 44784 38196 44790 38208
rect 51184 38196 51212 38372
rect 51810 38292 51816 38344
rect 51868 38332 51874 38344
rect 52733 38335 52791 38341
rect 52733 38332 52745 38335
rect 51868 38304 52745 38332
rect 51868 38292 51874 38304
rect 52733 38301 52745 38304
rect 52779 38301 52791 38335
rect 52733 38295 52791 38301
rect 51258 38224 51264 38276
rect 51316 38264 51322 38276
rect 52181 38267 52239 38273
rect 52181 38264 52193 38267
rect 51316 38236 52193 38264
rect 51316 38224 51322 38236
rect 52181 38233 52193 38236
rect 52227 38233 52239 38267
rect 52181 38227 52239 38233
rect 44784 38168 51212 38196
rect 51353 38199 51411 38205
rect 44784 38156 44790 38168
rect 51353 38165 51365 38199
rect 51399 38196 51411 38199
rect 51442 38196 51448 38208
rect 51399 38168 51448 38196
rect 51399 38165 51411 38168
rect 51353 38159 51411 38165
rect 51442 38156 51448 38168
rect 51500 38196 51506 38208
rect 52270 38196 52276 38208
rect 51500 38168 52276 38196
rect 51500 38156 51506 38168
rect 52270 38156 52276 38168
rect 52328 38156 52334 38208
rect 52840 38196 52868 38372
rect 52914 38292 52920 38344
rect 52972 38332 52978 38344
rect 53009 38335 53067 38341
rect 53009 38332 53021 38335
rect 52972 38304 53021 38332
rect 52972 38292 52978 38304
rect 53009 38301 53021 38304
rect 53055 38301 53067 38335
rect 53009 38295 53067 38301
rect 53116 38264 53144 38440
rect 53852 38440 53972 38468
rect 53374 38360 53380 38412
rect 53432 38400 53438 38412
rect 53852 38400 53880 38440
rect 54018 38428 54024 38480
rect 54076 38468 54082 38480
rect 54478 38468 54484 38480
rect 54076 38440 54484 38468
rect 54076 38428 54082 38440
rect 54478 38428 54484 38440
rect 54536 38428 54542 38480
rect 59262 38468 59268 38480
rect 59110 38440 59268 38468
rect 59262 38428 59268 38440
rect 59320 38428 59326 38480
rect 59538 38428 59544 38480
rect 59596 38428 59602 38480
rect 53432 38372 53880 38400
rect 53432 38360 53438 38372
rect 53926 38360 53932 38412
rect 53984 38400 53990 38412
rect 54389 38403 54447 38409
rect 54389 38400 54401 38403
rect 53984 38372 54401 38400
rect 53984 38360 53990 38372
rect 54389 38369 54401 38372
rect 54435 38369 54447 38403
rect 54389 38363 54447 38369
rect 55125 38403 55183 38409
rect 55125 38369 55137 38403
rect 55171 38400 55183 38403
rect 55214 38400 55220 38412
rect 55171 38372 55220 38400
rect 55171 38369 55183 38372
rect 55125 38363 55183 38369
rect 55214 38360 55220 38372
rect 55272 38360 55278 38412
rect 55766 38360 55772 38412
rect 55824 38360 55830 38412
rect 57425 38403 57483 38409
rect 57425 38369 57437 38403
rect 57471 38369 57483 38403
rect 64230 38400 64236 38412
rect 57425 38363 57483 38369
rect 59832 38372 64236 38400
rect 53193 38335 53251 38341
rect 53193 38301 53205 38335
rect 53239 38332 53251 38335
rect 53239 38304 54064 38332
rect 53239 38301 53251 38304
rect 53193 38295 53251 38301
rect 54036 38273 54064 38304
rect 54662 38292 54668 38344
rect 54720 38292 54726 38344
rect 56870 38292 56876 38344
rect 56928 38292 56934 38344
rect 57146 38292 57152 38344
rect 57204 38332 57210 38344
rect 57440 38332 57468 38363
rect 57204 38304 57468 38332
rect 57204 38292 57210 38304
rect 54021 38267 54079 38273
rect 53116 38236 53972 38264
rect 53374 38196 53380 38208
rect 52840 38168 53380 38196
rect 53374 38156 53380 38168
rect 53432 38156 53438 38208
rect 53834 38156 53840 38208
rect 53892 38156 53898 38208
rect 53944 38196 53972 38236
rect 54021 38233 54033 38267
rect 54067 38233 54079 38267
rect 57440 38264 57468 38304
rect 57698 38292 57704 38344
rect 57756 38332 57762 38344
rect 59832 38341 59860 38372
rect 64230 38360 64236 38372
rect 64288 38360 64294 38412
rect 57793 38335 57851 38341
rect 57793 38332 57805 38335
rect 57756 38304 57805 38332
rect 57756 38292 57762 38304
rect 57793 38301 57805 38304
rect 57839 38301 57851 38335
rect 59817 38335 59875 38341
rect 59817 38332 59829 38335
rect 57793 38295 57851 38301
rect 57900 38304 59829 38332
rect 57900 38264 57928 38304
rect 59817 38301 59829 38304
rect 59863 38301 59875 38335
rect 59817 38295 59875 38301
rect 60366 38292 60372 38344
rect 60424 38292 60430 38344
rect 60550 38292 60556 38344
rect 60608 38292 60614 38344
rect 60274 38264 60280 38276
rect 57440 38236 57928 38264
rect 59832 38236 60280 38264
rect 54021 38227 54079 38233
rect 57698 38196 57704 38208
rect 53944 38168 57704 38196
rect 57698 38156 57704 38168
rect 57756 38196 57762 38208
rect 59170 38196 59176 38208
rect 57756 38168 59176 38196
rect 57756 38156 57762 38168
rect 59170 38156 59176 38168
rect 59228 38196 59234 38208
rect 59832 38196 59860 38236
rect 60274 38224 60280 38236
rect 60332 38224 60338 38276
rect 59228 38168 59860 38196
rect 59228 38156 59234 38168
rect 59906 38156 59912 38208
rect 59964 38156 59970 38208
rect 59998 38156 60004 38208
rect 60056 38196 60062 38208
rect 63126 38196 63132 38208
rect 60056 38168 63132 38196
rect 60056 38156 60062 38168
rect 63126 38156 63132 38168
rect 63184 38156 63190 38208
rect 552 38106 66424 38128
rect 552 38054 1998 38106
rect 2050 38054 2062 38106
rect 2114 38054 2126 38106
rect 2178 38054 2190 38106
rect 2242 38054 2254 38106
rect 2306 38054 49998 38106
rect 50050 38054 50062 38106
rect 50114 38054 50126 38106
rect 50178 38054 50190 38106
rect 50242 38054 50254 38106
rect 50306 38054 66424 38106
rect 552 38032 66424 38054
rect 7466 37952 7472 38004
rect 7524 37952 7530 38004
rect 9306 37992 9312 38004
rect 8312 37964 9312 37992
rect 8113 37859 8171 37865
rect 8113 37825 8125 37859
rect 8159 37856 8171 37859
rect 8312 37856 8340 37964
rect 9306 37952 9312 37964
rect 9364 37952 9370 38004
rect 9674 37952 9680 38004
rect 9732 37992 9738 38004
rect 11514 37992 11520 38004
rect 9732 37964 11520 37992
rect 9732 37952 9738 37964
rect 8159 37828 8340 37856
rect 8389 37859 8447 37865
rect 8159 37825 8171 37828
rect 8113 37819 8171 37825
rect 8389 37825 8401 37859
rect 8435 37856 8447 37859
rect 8754 37856 8760 37868
rect 8435 37828 8760 37856
rect 8435 37825 8447 37828
rect 8389 37819 8447 37825
rect 8754 37816 8760 37828
rect 8812 37816 8818 37868
rect 10428 37865 10456 37964
rect 11514 37952 11520 37964
rect 11572 37992 11578 38004
rect 17221 37995 17279 38001
rect 11572 37964 17172 37992
rect 11572 37952 11578 37964
rect 14366 37884 14372 37936
rect 14424 37924 14430 37936
rect 14424 37896 14688 37924
rect 14424 37884 14430 37896
rect 10413 37859 10471 37865
rect 10413 37825 10425 37859
rect 10459 37825 10471 37859
rect 10413 37819 10471 37825
rect 10686 37816 10692 37868
rect 10744 37816 10750 37868
rect 10962 37816 10968 37868
rect 11020 37816 11026 37868
rect 13722 37816 13728 37868
rect 13780 37856 13786 37868
rect 13780 37828 14412 37856
rect 13780 37816 13786 37828
rect 7558 37748 7564 37800
rect 7616 37788 7622 37800
rect 7837 37791 7895 37797
rect 7837 37788 7849 37791
rect 7616 37760 7849 37788
rect 7616 37748 7622 37760
rect 7837 37757 7849 37760
rect 7883 37757 7895 37791
rect 12250 37788 12256 37800
rect 12098 37774 12256 37788
rect 7837 37751 7895 37757
rect 12084 37760 12256 37774
rect 8662 37680 8668 37732
rect 8720 37680 8726 37732
rect 9950 37720 9956 37732
rect 9890 37692 9956 37720
rect 9950 37680 9956 37692
rect 10008 37720 10014 37732
rect 10008 37692 11376 37720
rect 10008 37680 10014 37692
rect 7929 37655 7987 37661
rect 7929 37621 7941 37655
rect 7975 37652 7987 37655
rect 10962 37652 10968 37664
rect 7975 37624 10968 37652
rect 7975 37621 7987 37624
rect 7929 37615 7987 37621
rect 10962 37612 10968 37624
rect 11020 37612 11026 37664
rect 11348 37652 11376 37692
rect 12084 37652 12112 37760
rect 12250 37748 12256 37760
rect 12308 37788 12314 37800
rect 12308 37760 13676 37788
rect 12308 37748 12314 37760
rect 12618 37680 12624 37732
rect 12676 37720 12682 37732
rect 12713 37723 12771 37729
rect 12713 37720 12725 37723
rect 12676 37692 12725 37720
rect 12676 37680 12682 37692
rect 12713 37689 12725 37692
rect 12759 37689 12771 37723
rect 13648 37720 13676 37760
rect 14274 37720 14280 37732
rect 13648 37692 14280 37720
rect 12713 37683 12771 37689
rect 14274 37680 14280 37692
rect 14332 37680 14338 37732
rect 14384 37720 14412 37828
rect 14550 37816 14556 37868
rect 14608 37816 14614 37868
rect 14660 37865 14688 37896
rect 16482 37884 16488 37936
rect 16540 37924 16546 37936
rect 16669 37927 16727 37933
rect 16669 37924 16681 37927
rect 16540 37896 16681 37924
rect 16540 37884 16546 37896
rect 16669 37893 16681 37896
rect 16715 37924 16727 37927
rect 17144 37924 17172 37964
rect 17221 37961 17233 37995
rect 17267 37992 17279 37995
rect 17586 37992 17592 38004
rect 17267 37964 17592 37992
rect 17267 37961 17279 37964
rect 17221 37955 17279 37961
rect 17586 37952 17592 37964
rect 17644 37952 17650 38004
rect 18138 37952 18144 38004
rect 18196 37992 18202 38004
rect 18693 37995 18751 38001
rect 18693 37992 18705 37995
rect 18196 37964 18705 37992
rect 18196 37952 18202 37964
rect 18693 37961 18705 37964
rect 18739 37961 18751 37995
rect 18693 37955 18751 37961
rect 18782 37952 18788 38004
rect 18840 37992 18846 38004
rect 19334 37992 19340 38004
rect 18840 37964 19340 37992
rect 18840 37952 18846 37964
rect 19334 37952 19340 37964
rect 19392 37952 19398 38004
rect 19610 37952 19616 38004
rect 19668 37992 19674 38004
rect 19797 37995 19855 38001
rect 19797 37992 19809 37995
rect 19668 37964 19809 37992
rect 19668 37952 19674 37964
rect 19797 37961 19809 37964
rect 19843 37961 19855 37995
rect 20622 37992 20628 38004
rect 19797 37955 19855 37961
rect 19904 37964 20628 37992
rect 17770 37924 17776 37936
rect 16715 37896 17080 37924
rect 17144 37896 17776 37924
rect 16715 37893 16727 37896
rect 16669 37887 16727 37893
rect 14645 37859 14703 37865
rect 14645 37825 14657 37859
rect 14691 37825 14703 37859
rect 14645 37819 14703 37825
rect 14826 37816 14832 37868
rect 14884 37856 14890 37868
rect 14921 37859 14979 37865
rect 14921 37856 14933 37859
rect 14884 37828 14933 37856
rect 14884 37816 14890 37828
rect 14921 37825 14933 37828
rect 14967 37825 14979 37859
rect 14921 37819 14979 37825
rect 15194 37816 15200 37868
rect 15252 37816 15258 37868
rect 17052 37856 17080 37896
rect 17770 37884 17776 37896
rect 17828 37884 17834 37936
rect 17862 37884 17868 37936
rect 17920 37924 17926 37936
rect 19904 37924 19932 37964
rect 20622 37952 20628 37964
rect 20680 37952 20686 38004
rect 20714 37952 20720 38004
rect 20772 37952 20778 38004
rect 20990 37952 20996 38004
rect 21048 37992 21054 38004
rect 21048 37964 22094 37992
rect 21048 37952 21054 37964
rect 20732 37924 20760 37952
rect 17920 37896 19932 37924
rect 20456 37896 20760 37924
rect 22066 37924 22094 37964
rect 23566 37952 23572 38004
rect 23624 37992 23630 38004
rect 23845 37995 23903 38001
rect 23845 37992 23857 37995
rect 23624 37964 23857 37992
rect 23624 37952 23630 37964
rect 23845 37961 23857 37964
rect 23891 37961 23903 37995
rect 26326 37992 26332 38004
rect 23845 37955 23903 37961
rect 23952 37964 26332 37992
rect 23952 37924 23980 37964
rect 26326 37952 26332 37964
rect 26384 37952 26390 38004
rect 26510 37952 26516 38004
rect 26568 37952 26574 38004
rect 27798 37952 27804 38004
rect 27856 37992 27862 38004
rect 32030 37992 32036 38004
rect 27856 37964 32036 37992
rect 27856 37952 27862 37964
rect 32030 37952 32036 37964
rect 32088 37952 32094 38004
rect 33686 37992 33692 38004
rect 32140 37964 33692 37992
rect 26528 37924 26556 37952
rect 22066 37896 23980 37924
rect 26160 37896 26556 37924
rect 17920 37884 17926 37896
rect 20456 37865 20484 37896
rect 19337 37859 19395 37865
rect 17052 37828 19196 37856
rect 18138 37788 18144 37800
rect 16330 37760 18144 37788
rect 18138 37748 18144 37760
rect 18196 37748 18202 37800
rect 18506 37748 18512 37800
rect 18564 37748 18570 37800
rect 14384 37692 15516 37720
rect 11348 37624 12112 37652
rect 14090 37612 14096 37664
rect 14148 37612 14154 37664
rect 14461 37655 14519 37661
rect 14461 37621 14473 37655
rect 14507 37652 14519 37655
rect 15378 37652 15384 37664
rect 14507 37624 15384 37652
rect 14507 37621 14519 37624
rect 14461 37615 14519 37621
rect 15378 37612 15384 37624
rect 15436 37612 15442 37664
rect 15488 37652 15516 37692
rect 18782 37652 18788 37664
rect 15488 37624 18788 37652
rect 18782 37612 18788 37624
rect 18840 37612 18846 37664
rect 19058 37612 19064 37664
rect 19116 37612 19122 37664
rect 19168 37661 19196 37828
rect 19337 37825 19349 37859
rect 19383 37825 19395 37859
rect 19337 37819 19395 37825
rect 20441 37859 20499 37865
rect 20441 37825 20453 37859
rect 20487 37825 20499 37859
rect 20441 37819 20499 37825
rect 20625 37859 20683 37865
rect 20625 37825 20637 37859
rect 20671 37856 20683 37859
rect 24489 37859 24547 37865
rect 20671 37828 23428 37856
rect 20671 37825 20683 37828
rect 20625 37819 20683 37825
rect 19352 37720 19380 37819
rect 23400 37800 23428 37828
rect 24489 37825 24501 37859
rect 24535 37856 24547 37859
rect 26160 37856 26188 37896
rect 28258 37884 28264 37936
rect 28316 37884 28322 37936
rect 28902 37884 28908 37936
rect 28960 37924 28966 37936
rect 28997 37927 29055 37933
rect 28997 37924 29009 37927
rect 28960 37896 29009 37924
rect 28960 37884 28966 37896
rect 28997 37893 29009 37896
rect 29043 37893 29055 37927
rect 28997 37887 29055 37893
rect 31202 37884 31208 37936
rect 31260 37924 31266 37936
rect 32140 37924 32168 37964
rect 33686 37952 33692 37964
rect 33744 37952 33750 38004
rect 33781 37995 33839 38001
rect 33781 37961 33793 37995
rect 33827 37992 33839 37995
rect 33962 37992 33968 38004
rect 33827 37964 33968 37992
rect 33827 37961 33839 37964
rect 33781 37955 33839 37961
rect 33962 37952 33968 37964
rect 34020 37952 34026 38004
rect 36262 37992 36268 38004
rect 34164 37964 36268 37992
rect 34164 37924 34192 37964
rect 36262 37952 36268 37964
rect 36320 37952 36326 38004
rect 36906 37952 36912 38004
rect 36964 37952 36970 38004
rect 36998 37952 37004 38004
rect 37056 37992 37062 38004
rect 37056 37964 41000 37992
rect 37056 37952 37062 37964
rect 35069 37927 35127 37933
rect 35069 37924 35081 37927
rect 31260 37896 32168 37924
rect 33796 37896 34192 37924
rect 34256 37896 35081 37924
rect 31260 37884 31266 37896
rect 33796 37868 33824 37896
rect 34256 37868 34284 37896
rect 35069 37893 35081 37896
rect 35115 37893 35127 37927
rect 35069 37887 35127 37893
rect 36446 37884 36452 37936
rect 36504 37924 36510 37936
rect 40972 37924 41000 37964
rect 41230 37952 41236 38004
rect 41288 37952 41294 38004
rect 42702 37952 42708 38004
rect 42760 37992 42766 38004
rect 42797 37995 42855 38001
rect 42797 37992 42809 37995
rect 42760 37964 42809 37992
rect 42760 37952 42766 37964
rect 42797 37961 42809 37964
rect 42843 37961 42855 37995
rect 42797 37955 42855 37961
rect 43438 37952 43444 38004
rect 43496 37992 43502 38004
rect 43625 37995 43683 38001
rect 43625 37992 43637 37995
rect 43496 37964 43637 37992
rect 43496 37952 43502 37964
rect 43625 37961 43637 37964
rect 43671 37961 43683 37995
rect 43625 37955 43683 37961
rect 44542 37952 44548 38004
rect 44600 37952 44606 38004
rect 50798 37992 50804 38004
rect 45020 37964 50804 37992
rect 45020 37924 45048 37964
rect 50798 37952 50804 37964
rect 50856 37952 50862 38004
rect 51810 37952 51816 38004
rect 51868 37952 51874 38004
rect 57146 37992 57152 38004
rect 54588 37964 57152 37992
rect 36504 37896 40908 37924
rect 40972 37896 45048 37924
rect 46216 37896 47164 37924
rect 36504 37884 36510 37896
rect 24535 37828 26188 37856
rect 24535 37825 24547 37828
rect 24489 37819 24547 37825
rect 26234 37816 26240 37868
rect 26292 37856 26298 37868
rect 26513 37859 26571 37865
rect 26513 37856 26525 37859
rect 26292 37828 26525 37856
rect 26292 37816 26298 37828
rect 26513 37825 26525 37828
rect 26559 37825 26571 37859
rect 26513 37819 26571 37825
rect 26786 37816 26792 37868
rect 26844 37816 26850 37868
rect 27154 37816 27160 37868
rect 27212 37856 27218 37868
rect 29917 37859 29975 37865
rect 29917 37856 29929 37859
rect 27212 37828 29929 37856
rect 27212 37816 27218 37828
rect 29917 37825 29929 37828
rect 29963 37825 29975 37859
rect 29917 37819 29975 37825
rect 31386 37816 31392 37868
rect 31444 37816 31450 37868
rect 31754 37816 31760 37868
rect 31812 37856 31818 37868
rect 32022 37859 32080 37865
rect 32022 37856 32034 37859
rect 31812 37828 32034 37856
rect 31812 37816 31818 37828
rect 32022 37825 32034 37828
rect 32068 37825 32080 37859
rect 32022 37819 32080 37825
rect 32306 37816 32312 37868
rect 32364 37856 32370 37868
rect 32364 37828 33548 37856
rect 32364 37816 32370 37828
rect 20162 37748 20168 37800
rect 20220 37748 20226 37800
rect 23382 37748 23388 37800
rect 23440 37788 23446 37800
rect 24673 37791 24731 37797
rect 24673 37788 24685 37791
rect 23440 37760 24685 37788
rect 23440 37748 23446 37760
rect 24673 37757 24685 37760
rect 24719 37757 24731 37791
rect 24673 37751 24731 37757
rect 28258 37748 28264 37800
rect 28316 37788 28322 37800
rect 29549 37791 29607 37797
rect 29549 37788 29561 37791
rect 28316 37760 29561 37788
rect 28316 37748 28322 37760
rect 29549 37757 29561 37760
rect 29595 37757 29607 37791
rect 29549 37751 29607 37757
rect 20806 37720 20812 37732
rect 19352 37692 20812 37720
rect 20806 37680 20812 37692
rect 20864 37680 20870 37732
rect 20898 37680 20904 37732
rect 20956 37680 20962 37732
rect 21358 37680 21364 37732
rect 21416 37680 21422 37732
rect 22388 37692 24348 37720
rect 19153 37655 19211 37661
rect 19153 37621 19165 37655
rect 19199 37652 19211 37655
rect 19334 37652 19340 37664
rect 19199 37624 19340 37652
rect 19199 37621 19211 37624
rect 19153 37615 19211 37621
rect 19334 37612 19340 37624
rect 19392 37612 19398 37664
rect 20254 37612 20260 37664
rect 20312 37612 20318 37664
rect 21726 37612 21732 37664
rect 21784 37652 21790 37664
rect 22388 37661 22416 37692
rect 22373 37655 22431 37661
rect 22373 37652 22385 37655
rect 21784 37624 22385 37652
rect 21784 37612 21790 37624
rect 22373 37621 22385 37624
rect 22419 37621 22431 37655
rect 22373 37615 22431 37621
rect 24210 37612 24216 37664
rect 24268 37612 24274 37664
rect 24320 37661 24348 37692
rect 24946 37680 24952 37732
rect 25004 37680 25010 37732
rect 25038 37680 25044 37732
rect 25096 37720 25102 37732
rect 25096 37692 25438 37720
rect 25096 37680 25102 37692
rect 26326 37680 26332 37732
rect 26384 37720 26390 37732
rect 26384 37692 27278 37720
rect 26384 37680 26390 37692
rect 24305 37655 24363 37661
rect 24305 37621 24317 37655
rect 24351 37652 24363 37655
rect 24854 37652 24860 37664
rect 24351 37624 24860 37652
rect 24351 37621 24363 37624
rect 24305 37615 24363 37621
rect 24854 37612 24860 37624
rect 24912 37612 24918 37664
rect 26418 37612 26424 37664
rect 26476 37612 26482 37664
rect 27172 37652 27200 37692
rect 28074 37680 28080 37732
rect 28132 37720 28138 37732
rect 28132 37692 28994 37720
rect 28132 37680 28138 37692
rect 28442 37652 28448 37664
rect 27172 37624 28448 37652
rect 28442 37612 28448 37624
rect 28500 37612 28506 37664
rect 28966 37652 28994 37692
rect 30190 37680 30196 37732
rect 30248 37680 30254 37732
rect 31404 37720 31432 37816
rect 32214 37720 32220 37732
rect 31404 37706 32220 37720
rect 31418 37692 32220 37706
rect 32214 37680 32220 37692
rect 32272 37680 32278 37732
rect 32309 37723 32367 37729
rect 32309 37689 32321 37723
rect 32355 37720 32367 37723
rect 32398 37720 32404 37732
rect 32355 37692 32404 37720
rect 32355 37689 32367 37692
rect 32309 37683 32367 37689
rect 32398 37680 32404 37692
rect 32456 37680 32462 37732
rect 33520 37720 33548 37828
rect 33778 37816 33784 37868
rect 33836 37816 33842 37868
rect 34238 37816 34244 37868
rect 34296 37816 34302 37868
rect 34425 37859 34483 37865
rect 34425 37825 34437 37859
rect 34471 37856 34483 37859
rect 34698 37856 34704 37868
rect 34471 37828 34704 37856
rect 34471 37825 34483 37828
rect 34425 37819 34483 37825
rect 34698 37816 34704 37828
rect 34756 37816 34762 37868
rect 34974 37816 34980 37868
rect 35032 37856 35038 37868
rect 35158 37856 35164 37868
rect 35032 37828 35164 37856
rect 35032 37816 35038 37828
rect 35158 37816 35164 37828
rect 35216 37816 35222 37868
rect 35526 37816 35532 37868
rect 35584 37856 35590 37868
rect 38197 37859 38255 37865
rect 38197 37856 38209 37859
rect 35584 37828 38209 37856
rect 35584 37816 35590 37828
rect 38197 37825 38209 37828
rect 38243 37825 38255 37859
rect 38197 37819 38255 37825
rect 38565 37859 38623 37865
rect 38565 37825 38577 37859
rect 38611 37856 38623 37859
rect 39482 37856 39488 37868
rect 38611 37828 39488 37856
rect 38611 37825 38623 37828
rect 38565 37819 38623 37825
rect 33962 37748 33968 37800
rect 34020 37788 34026 37800
rect 34517 37791 34575 37797
rect 34517 37788 34529 37791
rect 34020 37760 34529 37788
rect 34020 37748 34026 37760
rect 34517 37757 34529 37760
rect 34563 37757 34575 37791
rect 34517 37751 34575 37757
rect 34624 37760 35204 37788
rect 33870 37720 33876 37732
rect 33520 37706 33876 37720
rect 33534 37692 33876 37706
rect 33870 37680 33876 37692
rect 33928 37720 33934 37732
rect 34624 37720 34652 37760
rect 35176 37732 35204 37760
rect 35250 37748 35256 37800
rect 35308 37788 35314 37800
rect 35621 37791 35679 37797
rect 35621 37788 35633 37791
rect 35308 37760 35633 37788
rect 35308 37748 35314 37760
rect 35621 37757 35633 37760
rect 35667 37757 35679 37791
rect 35621 37751 35679 37757
rect 35894 37748 35900 37800
rect 35952 37788 35958 37800
rect 37734 37788 37740 37800
rect 35952 37760 37740 37788
rect 35952 37748 35958 37760
rect 37734 37748 37740 37760
rect 37792 37748 37798 37800
rect 33928 37692 34652 37720
rect 33928 37680 33934 37692
rect 35158 37680 35164 37732
rect 35216 37680 35222 37732
rect 35342 37680 35348 37732
rect 35400 37720 35406 37732
rect 36998 37720 37004 37732
rect 35400 37692 37004 37720
rect 35400 37680 35406 37692
rect 36998 37680 37004 37692
rect 37056 37680 37062 37732
rect 38212 37720 38240 37819
rect 39482 37816 39488 37828
rect 39540 37816 39546 37868
rect 39945 37859 40003 37865
rect 39945 37825 39957 37859
rect 39991 37856 40003 37859
rect 40770 37856 40776 37868
rect 39991 37828 40776 37856
rect 39991 37825 40003 37828
rect 39945 37819 40003 37825
rect 40770 37816 40776 37828
rect 40828 37816 40834 37868
rect 38286 37748 38292 37800
rect 38344 37788 38350 37800
rect 38657 37791 38715 37797
rect 38657 37788 38669 37791
rect 38344 37760 38669 37788
rect 38344 37748 38350 37760
rect 38657 37757 38669 37760
rect 38703 37757 38715 37791
rect 38657 37751 38715 37757
rect 39114 37748 39120 37800
rect 39172 37788 39178 37800
rect 39669 37791 39727 37797
rect 39669 37788 39681 37791
rect 39172 37760 39681 37788
rect 39172 37748 39178 37760
rect 39669 37757 39681 37760
rect 39715 37757 39727 37791
rect 39669 37751 39727 37757
rect 39761 37791 39819 37797
rect 39761 37757 39773 37791
rect 39807 37788 39819 37791
rect 40126 37788 40132 37800
rect 39807 37760 40132 37788
rect 39807 37757 39819 37760
rect 39761 37751 39819 37757
rect 40126 37748 40132 37760
rect 40184 37748 40190 37800
rect 40494 37748 40500 37800
rect 40552 37788 40558 37800
rect 40552 37760 40816 37788
rect 40552 37748 40558 37760
rect 38749 37723 38807 37729
rect 38749 37720 38761 37723
rect 38212 37692 38761 37720
rect 38749 37689 38761 37692
rect 38795 37689 38807 37723
rect 40589 37723 40647 37729
rect 40589 37720 40601 37723
rect 38749 37683 38807 37689
rect 39132 37692 40601 37720
rect 31202 37652 31208 37664
rect 28966 37624 31208 37652
rect 31202 37612 31208 37624
rect 31260 37612 31266 37664
rect 31662 37612 31668 37664
rect 31720 37612 31726 37664
rect 32030 37612 32036 37664
rect 32088 37652 32094 37664
rect 34698 37652 34704 37664
rect 32088 37624 34704 37652
rect 32088 37612 32094 37624
rect 34698 37612 34704 37624
rect 34756 37612 34762 37664
rect 34882 37612 34888 37664
rect 34940 37612 34946 37664
rect 36170 37612 36176 37664
rect 36228 37652 36234 37664
rect 37274 37652 37280 37664
rect 36228 37624 37280 37652
rect 36228 37612 36234 37624
rect 37274 37612 37280 37624
rect 37332 37612 37338 37664
rect 39132 37661 39160 37692
rect 40589 37689 40601 37692
rect 40635 37689 40647 37723
rect 40589 37683 40647 37689
rect 39117 37655 39175 37661
rect 39117 37621 39129 37655
rect 39163 37621 39175 37655
rect 39117 37615 39175 37621
rect 39298 37612 39304 37664
rect 39356 37612 39362 37664
rect 40126 37612 40132 37664
rect 40184 37612 40190 37664
rect 40788 37652 40816 37760
rect 40880 37720 40908 37896
rect 42245 37859 42303 37865
rect 42245 37856 42257 37859
rect 41386 37828 42257 37856
rect 40954 37748 40960 37800
rect 41012 37788 41018 37800
rect 41386 37788 41414 37828
rect 42245 37825 42257 37828
rect 42291 37856 42303 37859
rect 42794 37856 42800 37868
rect 42291 37828 42800 37856
rect 42291 37825 42303 37828
rect 42245 37819 42303 37825
rect 42794 37816 42800 37828
rect 42852 37816 42858 37868
rect 43073 37859 43131 37865
rect 43073 37825 43085 37859
rect 43119 37856 43131 37859
rect 43346 37856 43352 37868
rect 43119 37828 43352 37856
rect 43119 37825 43131 37828
rect 43073 37819 43131 37825
rect 43346 37816 43352 37828
rect 43404 37816 43410 37868
rect 45278 37816 45284 37868
rect 45336 37856 45342 37868
rect 46216 37856 46244 37896
rect 45336 37828 46244 37856
rect 45336 37816 45342 37828
rect 41012 37760 41414 37788
rect 41012 37748 41018 37760
rect 41506 37748 41512 37800
rect 41564 37788 41570 37800
rect 41785 37791 41843 37797
rect 41785 37788 41797 37791
rect 41564 37760 41797 37788
rect 41564 37748 41570 37760
rect 41785 37757 41797 37760
rect 41831 37757 41843 37791
rect 41785 37751 41843 37757
rect 41966 37748 41972 37800
rect 42024 37788 42030 37800
rect 42429 37791 42487 37797
rect 42429 37788 42441 37791
rect 42024 37760 42441 37788
rect 42024 37748 42030 37760
rect 42429 37757 42441 37760
rect 42475 37788 42487 37791
rect 42702 37788 42708 37800
rect 42475 37760 42708 37788
rect 42475 37757 42487 37760
rect 42429 37751 42487 37757
rect 42702 37748 42708 37760
rect 42760 37788 42766 37800
rect 43165 37791 43223 37797
rect 43165 37788 43177 37791
rect 42760 37760 43177 37788
rect 42760 37748 42766 37760
rect 43165 37757 43177 37760
rect 43211 37757 43223 37791
rect 43165 37751 43223 37757
rect 43254 37748 43260 37800
rect 43312 37748 43318 37800
rect 46293 37791 46351 37797
rect 46293 37757 46305 37791
rect 46339 37788 46351 37791
rect 46934 37788 46940 37800
rect 46339 37760 46940 37788
rect 46339 37757 46351 37760
rect 46293 37751 46351 37757
rect 46934 37748 46940 37760
rect 46992 37748 46998 37800
rect 47136 37788 47164 37896
rect 48314 37856 48320 37868
rect 47412 37828 48320 37856
rect 47412 37788 47440 37828
rect 48314 37816 48320 37828
rect 48372 37816 48378 37868
rect 48406 37816 48412 37868
rect 48464 37816 48470 37868
rect 50065 37859 50123 37865
rect 50065 37825 50077 37859
rect 50111 37856 50123 37859
rect 51350 37856 51356 37868
rect 50111 37828 51356 37856
rect 50111 37825 50123 37828
rect 50065 37819 50123 37825
rect 47136 37760 47440 37788
rect 48678 37791 48736 37797
rect 48678 37757 48690 37791
rect 48724 37757 48736 37791
rect 48678 37751 48736 37757
rect 40880 37692 44772 37720
rect 41598 37652 41604 37664
rect 40788 37624 41604 37652
rect 41598 37612 41604 37624
rect 41656 37612 41662 37664
rect 42150 37612 42156 37664
rect 42208 37652 42214 37664
rect 42337 37655 42395 37661
rect 42337 37652 42349 37655
rect 42208 37624 42349 37652
rect 42208 37612 42214 37624
rect 42337 37621 42349 37624
rect 42383 37621 42395 37655
rect 44744 37652 44772 37692
rect 45278 37680 45284 37732
rect 45336 37680 45342 37732
rect 46014 37680 46020 37732
rect 46072 37680 46078 37732
rect 48314 37720 48320 37732
rect 46124 37692 47072 37720
rect 46124 37652 46152 37692
rect 44744 37624 46152 37652
rect 42337 37615 42395 37621
rect 46934 37612 46940 37664
rect 46992 37612 46998 37664
rect 47044 37652 47072 37692
rect 48056 37692 48320 37720
rect 48056 37652 48084 37692
rect 48314 37680 48320 37692
rect 48372 37680 48378 37732
rect 48700 37720 48728 37751
rect 49326 37748 49332 37800
rect 49384 37748 49390 37800
rect 50080 37720 50108 37819
rect 51350 37816 51356 37828
rect 51408 37816 51414 37868
rect 54588 37865 54616 37964
rect 57146 37952 57152 37964
rect 57204 37952 57210 38004
rect 57790 37952 57796 38004
rect 57848 37952 57854 38004
rect 57900 37964 60136 37992
rect 55950 37884 55956 37936
rect 56008 37924 56014 37936
rect 56045 37927 56103 37933
rect 56045 37924 56057 37927
rect 56008 37896 56057 37924
rect 56008 37884 56014 37896
rect 56045 37893 56057 37896
rect 56091 37893 56103 37927
rect 56045 37887 56103 37893
rect 56152 37896 56364 37924
rect 54573 37859 54631 37865
rect 54573 37825 54585 37859
rect 54619 37825 54631 37859
rect 54573 37819 54631 37825
rect 54662 37816 54668 37868
rect 54720 37856 54726 37868
rect 55493 37859 55551 37865
rect 55493 37856 55505 37859
rect 54720 37828 55505 37856
rect 54720 37816 54726 37828
rect 55493 37825 55505 37828
rect 55539 37856 55551 37859
rect 56152 37856 56180 37896
rect 55539 37828 56180 37856
rect 55539 37825 55551 37828
rect 55493 37819 55551 37825
rect 56226 37816 56232 37868
rect 56284 37816 56290 37868
rect 56336 37856 56364 37896
rect 56870 37884 56876 37936
rect 56928 37884 56934 37936
rect 57241 37859 57299 37865
rect 57241 37856 57253 37859
rect 56336 37828 57253 37856
rect 57241 37825 57253 37828
rect 57287 37856 57299 37859
rect 57900 37856 57928 37964
rect 57287 37828 57928 37856
rect 57287 37825 57299 37828
rect 57241 37819 57299 37825
rect 58158 37816 58164 37868
rect 58216 37816 58222 37868
rect 58250 37816 58256 37868
rect 58308 37856 58314 37868
rect 60108 37865 60136 37964
rect 60366 37952 60372 38004
rect 60424 37992 60430 38004
rect 60645 37995 60703 38001
rect 60645 37992 60657 37995
rect 60424 37964 60657 37992
rect 60424 37952 60430 37964
rect 60645 37961 60657 37964
rect 60691 37961 60703 37995
rect 60645 37955 60703 37961
rect 60093 37859 60151 37865
rect 58308 37828 59860 37856
rect 58308 37816 58314 37828
rect 53006 37788 53012 37800
rect 51474 37760 53012 37788
rect 53006 37748 53012 37760
rect 53064 37788 53070 37800
rect 53064 37760 53222 37788
rect 53064 37748 53070 37760
rect 55214 37748 55220 37800
rect 55272 37788 55278 37800
rect 55677 37791 55735 37797
rect 55677 37788 55689 37791
rect 55272 37760 55689 37788
rect 55272 37748 55278 37760
rect 55677 37757 55689 37760
rect 55723 37757 55735 37791
rect 55677 37751 55735 37757
rect 48700 37692 50108 37720
rect 50338 37680 50344 37732
rect 50396 37680 50402 37732
rect 52546 37680 52552 37732
rect 52604 37680 52610 37732
rect 54294 37680 54300 37732
rect 54352 37680 54358 37732
rect 55692 37720 55720 37751
rect 56042 37748 56048 37800
rect 56100 37788 56106 37800
rect 57885 37791 57943 37797
rect 57885 37788 57897 37791
rect 56100 37760 57897 37788
rect 56100 37748 56106 37760
rect 57885 37757 57897 37760
rect 57931 37757 57943 37791
rect 57885 37751 57943 37757
rect 59262 37748 59268 37800
rect 59320 37748 59326 37800
rect 56413 37723 56471 37729
rect 56413 37720 56425 37723
rect 55692 37692 56425 37720
rect 56413 37689 56425 37692
rect 56459 37689 56471 37723
rect 56413 37683 56471 37689
rect 56505 37723 56563 37729
rect 56505 37689 56517 37723
rect 56551 37720 56563 37723
rect 56778 37720 56784 37732
rect 56551 37692 56784 37720
rect 56551 37689 56563 37692
rect 56505 37683 56563 37689
rect 47044 37624 48084 37652
rect 48222 37612 48228 37664
rect 48280 37652 48286 37664
rect 48777 37655 48835 37661
rect 48777 37652 48789 37655
rect 48280 37624 48789 37652
rect 48280 37612 48286 37624
rect 48777 37621 48789 37624
rect 48823 37621 48835 37655
rect 48777 37615 48835 37621
rect 53650 37612 53656 37664
rect 53708 37652 53714 37664
rect 55585 37655 55643 37661
rect 55585 37652 55597 37655
rect 53708 37624 55597 37652
rect 53708 37612 53714 37624
rect 55585 37621 55597 37624
rect 55631 37621 55643 37655
rect 56428 37652 56456 37683
rect 56778 37680 56784 37692
rect 56836 37680 56842 37732
rect 56870 37680 56876 37732
rect 56928 37720 56934 37732
rect 57425 37723 57483 37729
rect 57425 37720 57437 37723
rect 56928 37692 57437 37720
rect 56928 37680 56934 37692
rect 57425 37689 57437 37692
rect 57471 37720 57483 37723
rect 58250 37720 58256 37732
rect 57471 37692 58256 37720
rect 57471 37689 57483 37692
rect 57425 37683 57483 37689
rect 58250 37680 58256 37692
rect 58308 37680 58314 37732
rect 59832 37664 59860 37828
rect 60093 37825 60105 37859
rect 60139 37856 60151 37859
rect 63954 37856 63960 37868
rect 60139 37828 63960 37856
rect 60139 37825 60151 37828
rect 60093 37819 60151 37825
rect 63954 37816 63960 37828
rect 64012 37816 64018 37868
rect 60274 37748 60280 37800
rect 60332 37748 60338 37800
rect 62482 37748 62488 37800
rect 62540 37788 62546 37800
rect 63402 37788 63408 37800
rect 62540 37760 63408 37788
rect 62540 37748 62546 37760
rect 63402 37748 63408 37760
rect 63460 37748 63466 37800
rect 57333 37655 57391 37661
rect 57333 37652 57345 37655
rect 56428 37624 57345 37652
rect 55585 37615 55643 37621
rect 57333 37621 57345 37624
rect 57379 37621 57391 37655
rect 57333 37615 57391 37621
rect 58066 37612 58072 37664
rect 58124 37652 58130 37664
rect 59630 37652 59636 37664
rect 58124 37624 59636 37652
rect 58124 37612 58130 37624
rect 59630 37612 59636 37624
rect 59688 37612 59694 37664
rect 59814 37612 59820 37664
rect 59872 37652 59878 37664
rect 60185 37655 60243 37661
rect 60185 37652 60197 37655
rect 59872 37624 60197 37652
rect 59872 37612 59878 37624
rect 60185 37621 60197 37624
rect 60231 37621 60243 37655
rect 60185 37615 60243 37621
rect 64046 37612 64052 37664
rect 64104 37612 64110 37664
rect 552 37562 66424 37584
rect 552 37510 2918 37562
rect 2970 37510 2982 37562
rect 3034 37510 3046 37562
rect 3098 37510 3110 37562
rect 3162 37510 3174 37562
rect 3226 37510 50918 37562
rect 50970 37510 50982 37562
rect 51034 37510 51046 37562
rect 51098 37510 51110 37562
rect 51162 37510 51174 37562
rect 51226 37510 65258 37562
rect 65310 37510 65322 37562
rect 65374 37510 65386 37562
rect 65438 37510 65450 37562
rect 65502 37510 65514 37562
rect 65566 37510 66424 37562
rect 552 37488 66424 37510
rect 8662 37408 8668 37460
rect 8720 37448 8726 37460
rect 9033 37451 9091 37457
rect 9033 37448 9045 37451
rect 8720 37420 9045 37448
rect 8720 37408 8726 37420
rect 9033 37417 9045 37420
rect 9079 37417 9091 37451
rect 9033 37411 9091 37417
rect 9493 37451 9551 37457
rect 9493 37417 9505 37451
rect 9539 37448 9551 37451
rect 9674 37448 9680 37460
rect 9539 37420 9680 37448
rect 9539 37417 9551 37420
rect 9493 37411 9551 37417
rect 9674 37408 9680 37420
rect 9732 37408 9738 37460
rect 10962 37408 10968 37460
rect 11020 37408 11026 37460
rect 11330 37408 11336 37460
rect 11388 37448 11394 37460
rect 12253 37451 12311 37457
rect 12253 37448 12265 37451
rect 11388 37420 12265 37448
rect 11388 37408 11394 37420
rect 12253 37417 12265 37420
rect 12299 37417 12311 37451
rect 12713 37451 12771 37457
rect 12713 37448 12725 37451
rect 12253 37411 12311 37417
rect 12406 37420 12725 37448
rect 12406 37392 12434 37420
rect 12713 37417 12725 37420
rect 12759 37448 12771 37451
rect 12759 37420 15240 37448
rect 12759 37417 12771 37420
rect 12713 37411 12771 37417
rect 8846 37340 8852 37392
rect 8904 37380 8910 37392
rect 9401 37383 9459 37389
rect 9401 37380 9413 37383
rect 8904 37352 9413 37380
rect 8904 37340 8910 37352
rect 9401 37349 9413 37352
rect 9447 37349 9459 37383
rect 11514 37380 11520 37392
rect 9401 37343 9459 37349
rect 11348 37352 11520 37380
rect 11348 37321 11376 37352
rect 11514 37340 11520 37352
rect 11572 37340 11578 37392
rect 12342 37340 12348 37392
rect 12400 37352 12434 37392
rect 12400 37340 12406 37352
rect 12618 37340 12624 37392
rect 12676 37340 12682 37392
rect 13817 37383 13875 37389
rect 13817 37349 13829 37383
rect 13863 37380 13875 37383
rect 14090 37380 14096 37392
rect 13863 37352 14096 37380
rect 13863 37349 13875 37352
rect 13817 37343 13875 37349
rect 14090 37340 14096 37352
rect 14148 37340 14154 37392
rect 14274 37340 14280 37392
rect 14332 37340 14338 37392
rect 15212 37380 15240 37420
rect 15286 37408 15292 37460
rect 15344 37408 15350 37460
rect 17678 37448 17684 37460
rect 15764 37420 17684 37448
rect 15764 37380 15792 37420
rect 17678 37408 17684 37420
rect 17736 37408 17742 37460
rect 18414 37408 18420 37460
rect 18472 37448 18478 37460
rect 19061 37451 19119 37457
rect 19061 37448 19073 37451
rect 18472 37420 19073 37448
rect 18472 37408 18478 37420
rect 19061 37417 19073 37420
rect 19107 37417 19119 37451
rect 19061 37411 19119 37417
rect 20254 37408 20260 37460
rect 20312 37448 20318 37460
rect 21361 37451 21419 37457
rect 21361 37448 21373 37451
rect 20312 37420 21373 37448
rect 20312 37408 20318 37420
rect 21361 37417 21373 37420
rect 21407 37417 21419 37451
rect 21361 37411 21419 37417
rect 21726 37408 21732 37460
rect 21784 37408 21790 37460
rect 24946 37408 24952 37460
rect 25004 37448 25010 37460
rect 25501 37451 25559 37457
rect 25501 37448 25513 37451
rect 25004 37420 25513 37448
rect 25004 37408 25010 37420
rect 25501 37417 25513 37420
rect 25547 37417 25559 37451
rect 25501 37411 25559 37417
rect 25866 37408 25872 37460
rect 25924 37408 25930 37460
rect 25958 37408 25964 37460
rect 26016 37408 26022 37460
rect 26142 37408 26148 37460
rect 26200 37448 26206 37460
rect 26421 37451 26479 37457
rect 26421 37448 26433 37451
rect 26200 37420 26433 37448
rect 26200 37408 26206 37420
rect 26421 37417 26433 37420
rect 26467 37417 26479 37451
rect 26421 37411 26479 37417
rect 26881 37451 26939 37457
rect 26881 37417 26893 37451
rect 26927 37448 26939 37451
rect 27430 37448 27436 37460
rect 26927 37420 27436 37448
rect 26927 37417 26939 37420
rect 26881 37411 26939 37417
rect 27430 37408 27436 37420
rect 27488 37408 27494 37460
rect 27706 37408 27712 37460
rect 27764 37448 27770 37460
rect 27893 37451 27951 37457
rect 27893 37448 27905 37451
rect 27764 37420 27905 37448
rect 27764 37408 27770 37420
rect 27893 37417 27905 37420
rect 27939 37417 27951 37451
rect 27893 37411 27951 37417
rect 28261 37451 28319 37457
rect 28261 37417 28273 37451
rect 28307 37448 28319 37451
rect 28902 37448 28908 37460
rect 28307 37420 28908 37448
rect 28307 37417 28319 37420
rect 28261 37411 28319 37417
rect 28902 37408 28908 37420
rect 28960 37408 28966 37460
rect 30190 37408 30196 37460
rect 30248 37448 30254 37460
rect 30377 37451 30435 37457
rect 30377 37448 30389 37451
rect 30248 37420 30389 37448
rect 30248 37408 30254 37420
rect 30377 37417 30389 37420
rect 30423 37417 30435 37451
rect 30377 37411 30435 37417
rect 30742 37408 30748 37460
rect 30800 37408 30806 37460
rect 30834 37408 30840 37460
rect 30892 37448 30898 37460
rect 32306 37448 32312 37460
rect 30892 37420 32312 37448
rect 30892 37408 30898 37420
rect 32306 37408 32312 37420
rect 32364 37408 32370 37460
rect 32398 37408 32404 37460
rect 32456 37408 32462 37460
rect 32861 37451 32919 37457
rect 32861 37417 32873 37451
rect 32907 37448 32919 37451
rect 33229 37451 33287 37457
rect 33229 37448 33241 37451
rect 32907 37420 33241 37448
rect 32907 37417 32919 37420
rect 32861 37411 32919 37417
rect 33229 37417 33241 37420
rect 33275 37417 33287 37451
rect 36446 37448 36452 37460
rect 33229 37411 33287 37417
rect 33428 37420 36452 37448
rect 15212 37352 15792 37380
rect 20714 37340 20720 37392
rect 20772 37380 20778 37392
rect 32769 37383 32827 37389
rect 20772 37352 32720 37380
rect 20772 37340 20778 37352
rect 11333 37315 11391 37321
rect 11333 37281 11345 37315
rect 11379 37281 11391 37315
rect 11333 37275 11391 37281
rect 11425 37315 11483 37321
rect 11425 37281 11437 37315
rect 11471 37312 11483 37315
rect 12636 37312 12664 37340
rect 11471 37284 12664 37312
rect 11471 37281 11483 37284
rect 11425 37275 11483 37281
rect 13538 37272 13544 37324
rect 13596 37272 13602 37324
rect 16758 37272 16764 37324
rect 16816 37272 16822 37324
rect 18138 37272 18144 37324
rect 18196 37272 18202 37324
rect 19058 37312 19064 37324
rect 18800 37284 19064 37312
rect 9582 37204 9588 37256
rect 9640 37204 9646 37256
rect 11238 37204 11244 37256
rect 11296 37244 11302 37256
rect 11517 37247 11575 37253
rect 11517 37244 11529 37247
rect 11296 37216 11529 37244
rect 11296 37204 11302 37216
rect 11517 37213 11529 37216
rect 11563 37244 11575 37247
rect 12805 37247 12863 37253
rect 12805 37244 12817 37247
rect 11563 37216 12817 37244
rect 11563 37213 11575 37216
rect 11517 37207 11575 37213
rect 12805 37213 12817 37216
rect 12851 37213 12863 37247
rect 12805 37207 12863 37213
rect 17037 37247 17095 37253
rect 17037 37213 17049 37247
rect 17083 37244 17095 37247
rect 17083 37216 18736 37244
rect 17083 37213 17095 37216
rect 17037 37207 17095 37213
rect 18708 37185 18736 37216
rect 18693 37179 18751 37185
rect 18693 37145 18705 37179
rect 18739 37145 18751 37179
rect 18693 37139 18751 37145
rect 18509 37111 18567 37117
rect 18509 37077 18521 37111
rect 18555 37108 18567 37111
rect 18800 37108 18828 37284
rect 19058 37272 19064 37284
rect 19116 37312 19122 37324
rect 19153 37315 19211 37321
rect 19153 37312 19165 37315
rect 19116 37284 19165 37312
rect 19116 37272 19122 37284
rect 19153 37281 19165 37284
rect 19199 37312 19211 37315
rect 21821 37315 21879 37321
rect 21821 37312 21833 37315
rect 19199 37284 21833 37312
rect 19199 37281 19211 37284
rect 19153 37275 19211 37281
rect 21821 37281 21833 37284
rect 21867 37312 21879 37315
rect 23198 37312 23204 37324
rect 21867 37284 23204 37312
rect 21867 37281 21879 37284
rect 21821 37275 21879 37281
rect 23198 37272 23204 37284
rect 23256 37272 23262 37324
rect 25038 37272 25044 37324
rect 25096 37312 25102 37324
rect 26326 37312 26332 37324
rect 25096 37284 26332 37312
rect 25096 37272 25102 37284
rect 26326 37272 26332 37284
rect 26384 37272 26390 37324
rect 26418 37272 26424 37324
rect 26476 37312 26482 37324
rect 26789 37315 26847 37321
rect 26789 37312 26801 37315
rect 26476 37284 26801 37312
rect 26476 37272 26482 37284
rect 26789 37281 26801 37284
rect 26835 37312 26847 37315
rect 28353 37315 28411 37321
rect 28353 37312 28365 37315
rect 26835 37284 28365 37312
rect 26835 37281 26847 37284
rect 26789 37275 26847 37281
rect 28353 37281 28365 37284
rect 28399 37312 28411 37315
rect 30742 37312 30748 37324
rect 28399 37284 30748 37312
rect 28399 37281 28411 37284
rect 28353 37275 28411 37281
rect 30742 37272 30748 37284
rect 30800 37272 30806 37324
rect 30837 37315 30895 37321
rect 30837 37281 30849 37315
rect 30883 37312 30895 37315
rect 31573 37315 31631 37321
rect 31573 37312 31585 37315
rect 30883 37284 31585 37312
rect 30883 37281 30895 37284
rect 30837 37275 30895 37281
rect 31573 37281 31585 37284
rect 31619 37281 31631 37315
rect 31573 37275 31631 37281
rect 31662 37272 31668 37324
rect 31720 37312 31726 37324
rect 32125 37315 32183 37321
rect 32125 37312 32137 37315
rect 31720 37284 32137 37312
rect 31720 37272 31726 37284
rect 32125 37281 32137 37284
rect 32171 37281 32183 37315
rect 32692 37312 32720 37352
rect 32769 37349 32781 37383
rect 32815 37380 32827 37383
rect 33318 37380 33324 37392
rect 32815 37352 33324 37380
rect 32815 37349 32827 37352
rect 32769 37343 32827 37349
rect 33318 37340 33324 37352
rect 33376 37340 33382 37392
rect 33428 37312 33456 37420
rect 36446 37408 36452 37420
rect 36504 37408 36510 37460
rect 36541 37451 36599 37457
rect 36541 37417 36553 37451
rect 36587 37448 36599 37451
rect 36814 37448 36820 37460
rect 36587 37420 36820 37448
rect 36587 37417 36599 37420
rect 36541 37411 36599 37417
rect 36814 37408 36820 37420
rect 36872 37408 36878 37460
rect 41690 37448 41696 37460
rect 39960 37420 41696 37448
rect 33502 37340 33508 37392
rect 33560 37380 33566 37392
rect 33689 37383 33747 37389
rect 33689 37380 33701 37383
rect 33560 37352 33701 37380
rect 33560 37340 33566 37352
rect 33689 37349 33701 37352
rect 33735 37349 33747 37383
rect 33689 37343 33747 37349
rect 34974 37340 34980 37392
rect 35032 37380 35038 37392
rect 35069 37383 35127 37389
rect 35069 37380 35081 37383
rect 35032 37352 35081 37380
rect 35032 37340 35038 37352
rect 35069 37349 35081 37352
rect 35115 37349 35127 37383
rect 35069 37343 35127 37349
rect 35158 37340 35164 37392
rect 35216 37380 35222 37392
rect 35216 37352 35558 37380
rect 35216 37340 35222 37352
rect 36722 37340 36728 37392
rect 36780 37340 36786 37392
rect 32692 37284 33456 37312
rect 32125 37275 32183 37281
rect 33594 37272 33600 37324
rect 33652 37272 33658 37324
rect 34790 37272 34796 37324
rect 34848 37272 34854 37324
rect 39960 37321 39988 37420
rect 41690 37408 41696 37420
rect 41748 37408 41754 37460
rect 42702 37408 42708 37460
rect 42760 37448 42766 37460
rect 44729 37451 44787 37457
rect 44729 37448 44741 37451
rect 42760 37420 44741 37448
rect 42760 37408 42766 37420
rect 44729 37417 44741 37420
rect 44775 37417 44787 37451
rect 44729 37411 44787 37417
rect 44910 37408 44916 37460
rect 44968 37448 44974 37460
rect 45189 37451 45247 37457
rect 45189 37448 45201 37451
rect 44968 37420 45201 37448
rect 44968 37408 44974 37420
rect 45189 37417 45201 37420
rect 45235 37417 45247 37451
rect 45189 37411 45247 37417
rect 45646 37408 45652 37460
rect 45704 37408 45710 37460
rect 46014 37408 46020 37460
rect 46072 37408 46078 37460
rect 47762 37408 47768 37460
rect 47820 37408 47826 37460
rect 48222 37408 48228 37460
rect 48280 37408 48286 37460
rect 48498 37408 48504 37460
rect 48556 37448 48562 37460
rect 48593 37451 48651 37457
rect 48593 37448 48605 37451
rect 48556 37420 48605 37448
rect 48556 37408 48562 37420
rect 48593 37417 48605 37420
rect 48639 37417 48651 37451
rect 48593 37411 48651 37417
rect 49973 37451 50031 37457
rect 49973 37417 49985 37451
rect 50019 37448 50031 37451
rect 50246 37448 50252 37460
rect 50019 37420 50252 37448
rect 50019 37417 50031 37420
rect 49973 37411 50031 37417
rect 50246 37408 50252 37420
rect 50304 37408 50310 37460
rect 50338 37408 50344 37460
rect 50396 37448 50402 37460
rect 50893 37451 50951 37457
rect 50893 37448 50905 37451
rect 50396 37420 50905 37448
rect 50396 37408 50402 37420
rect 50893 37417 50905 37420
rect 50939 37417 50951 37451
rect 50893 37411 50951 37417
rect 51258 37408 51264 37460
rect 51316 37408 51322 37460
rect 51353 37451 51411 37457
rect 51353 37417 51365 37451
rect 51399 37448 51411 37451
rect 52181 37451 52239 37457
rect 52181 37448 52193 37451
rect 51399 37420 52193 37448
rect 51399 37417 51411 37420
rect 51353 37411 51411 37417
rect 52181 37417 52193 37420
rect 52227 37417 52239 37451
rect 52181 37411 52239 37417
rect 52270 37408 52276 37460
rect 52328 37448 52334 37460
rect 52549 37451 52607 37457
rect 52549 37448 52561 37451
rect 52328 37420 52561 37448
rect 52328 37408 52334 37420
rect 52549 37417 52561 37420
rect 52595 37417 52607 37451
rect 52549 37411 52607 37417
rect 52730 37408 52736 37460
rect 52788 37448 52794 37460
rect 53190 37448 53196 37460
rect 52788 37420 53196 37448
rect 52788 37408 52794 37420
rect 53190 37408 53196 37420
rect 53248 37408 53254 37460
rect 53558 37408 53564 37460
rect 53616 37448 53622 37460
rect 53745 37451 53803 37457
rect 53745 37448 53757 37451
rect 53616 37420 53757 37448
rect 53616 37408 53622 37420
rect 53745 37417 53757 37420
rect 53791 37417 53803 37451
rect 53745 37411 53803 37417
rect 54113 37451 54171 37457
rect 54113 37417 54125 37451
rect 54159 37448 54171 37451
rect 54294 37448 54300 37460
rect 54159 37420 54300 37448
rect 54159 37417 54171 37420
rect 54113 37411 54171 37417
rect 54294 37408 54300 37420
rect 54352 37408 54358 37460
rect 56686 37408 56692 37460
rect 56744 37408 56750 37460
rect 56781 37451 56839 37457
rect 56781 37417 56793 37451
rect 56827 37448 56839 37451
rect 58066 37448 58072 37460
rect 56827 37420 58072 37448
rect 56827 37417 56839 37420
rect 56781 37411 56839 37417
rect 58066 37408 58072 37420
rect 58124 37408 58130 37460
rect 58176 37420 59216 37448
rect 40126 37340 40132 37392
rect 40184 37380 40190 37392
rect 40221 37383 40279 37389
rect 40221 37380 40233 37383
rect 40184 37352 40233 37380
rect 40184 37340 40190 37352
rect 40221 37349 40233 37352
rect 40267 37349 40279 37383
rect 40221 37343 40279 37349
rect 44082 37340 44088 37392
rect 44140 37380 44146 37392
rect 44140 37352 44956 37380
rect 44140 37340 44146 37352
rect 39945 37315 40003 37321
rect 39945 37281 39957 37315
rect 39991 37281 40003 37315
rect 39945 37275 40003 37281
rect 41230 37272 41236 37324
rect 41288 37272 41294 37324
rect 41322 37272 41328 37324
rect 41380 37272 41386 37324
rect 43346 37312 43352 37324
rect 41432 37284 43352 37312
rect 19242 37204 19248 37256
rect 19300 37204 19306 37256
rect 20806 37204 20812 37256
rect 20864 37244 20870 37256
rect 21913 37247 21971 37253
rect 21913 37244 21925 37247
rect 20864 37216 21925 37244
rect 20864 37204 20870 37216
rect 21913 37213 21925 37216
rect 21959 37213 21971 37247
rect 21913 37207 21971 37213
rect 26145 37247 26203 37253
rect 26145 37213 26157 37247
rect 26191 37213 26203 37247
rect 26145 37207 26203 37213
rect 20622 37136 20628 37188
rect 20680 37176 20686 37188
rect 25222 37176 25228 37188
rect 20680 37148 25228 37176
rect 20680 37136 20686 37148
rect 25222 37136 25228 37148
rect 25280 37136 25286 37188
rect 26160 37176 26188 37207
rect 26510 37204 26516 37256
rect 26568 37244 26574 37256
rect 27065 37247 27123 37253
rect 27065 37244 27077 37247
rect 26568 37216 27077 37244
rect 26568 37204 26574 37216
rect 27065 37213 27077 37216
rect 27111 37244 27123 37247
rect 28537 37247 28595 37253
rect 28537 37244 28549 37247
rect 27111 37216 28549 37244
rect 27111 37213 27123 37216
rect 27065 37207 27123 37213
rect 28537 37213 28549 37216
rect 28583 37244 28595 37247
rect 28718 37244 28724 37256
rect 28583 37216 28724 37244
rect 28583 37213 28595 37216
rect 28537 37207 28595 37213
rect 28718 37204 28724 37216
rect 28776 37204 28782 37256
rect 31021 37247 31079 37253
rect 31021 37213 31033 37247
rect 31067 37244 31079 37247
rect 31478 37244 31484 37256
rect 31067 37216 31484 37244
rect 31067 37213 31079 37216
rect 31021 37207 31079 37213
rect 31478 37204 31484 37216
rect 31536 37204 31542 37256
rect 33045 37247 33103 37253
rect 33045 37244 33057 37247
rect 31726 37216 33057 37244
rect 27522 37176 27528 37188
rect 26160 37148 27528 37176
rect 27522 37136 27528 37148
rect 27580 37136 27586 37188
rect 30282 37136 30288 37188
rect 30340 37176 30346 37188
rect 31726 37176 31754 37216
rect 33045 37213 33057 37216
rect 33091 37244 33103 37247
rect 33134 37244 33140 37256
rect 33091 37216 33140 37244
rect 33091 37213 33103 37216
rect 33045 37207 33103 37213
rect 33134 37204 33140 37216
rect 33192 37204 33198 37256
rect 33873 37247 33931 37253
rect 33873 37213 33885 37247
rect 33919 37244 33931 37247
rect 35066 37244 35072 37256
rect 33919 37216 35072 37244
rect 33919 37213 33931 37216
rect 33873 37207 33931 37213
rect 35066 37204 35072 37216
rect 35124 37244 35130 37256
rect 35710 37244 35716 37256
rect 35124 37216 35716 37244
rect 35124 37204 35130 37216
rect 35710 37204 35716 37216
rect 35768 37204 35774 37256
rect 38470 37204 38476 37256
rect 38528 37204 38534 37256
rect 41248 37244 41276 37272
rect 41432 37244 41460 37284
rect 43346 37272 43352 37284
rect 43404 37272 43410 37324
rect 44634 37272 44640 37324
rect 44692 37312 44698 37324
rect 44818 37312 44824 37324
rect 44692 37284 44824 37312
rect 44692 37272 44698 37284
rect 44818 37272 44824 37284
rect 44876 37272 44882 37324
rect 44928 37312 44956 37352
rect 45094 37340 45100 37392
rect 45152 37380 45158 37392
rect 45554 37380 45560 37392
rect 45152 37352 45560 37380
rect 45152 37340 45158 37352
rect 45554 37340 45560 37352
rect 45612 37340 45618 37392
rect 46934 37340 46940 37392
rect 46992 37380 46998 37392
rect 47305 37383 47363 37389
rect 47305 37380 47317 37383
rect 46992 37352 47317 37380
rect 46992 37340 46998 37352
rect 47305 37349 47317 37352
rect 47351 37380 47363 37383
rect 49326 37380 49332 37392
rect 47351 37352 49332 37380
rect 47351 37349 47363 37352
rect 47305 37343 47363 37349
rect 49326 37340 49332 37352
rect 49384 37340 49390 37392
rect 50433 37383 50491 37389
rect 50433 37349 50445 37383
rect 50479 37380 50491 37383
rect 51810 37380 51816 37392
rect 50479 37352 51816 37380
rect 50479 37349 50491 37352
rect 50433 37343 50491 37349
rect 51810 37340 51816 37352
rect 51868 37340 51874 37392
rect 52641 37383 52699 37389
rect 52641 37349 52653 37383
rect 52687 37380 52699 37383
rect 58176 37380 58204 37420
rect 52687 37352 58204 37380
rect 52687 37349 52699 37352
rect 52641 37343 52699 37349
rect 47397 37315 47455 37321
rect 47397 37312 47409 37315
rect 44928 37284 47409 37312
rect 47397 37281 47409 37284
rect 47443 37281 47455 37315
rect 49789 37315 49847 37321
rect 49789 37312 49801 37315
rect 47397 37275 47455 37281
rect 47504 37284 49801 37312
rect 41248 37216 41460 37244
rect 42794 37204 42800 37256
rect 42852 37244 42858 37256
rect 44545 37247 44603 37253
rect 44545 37244 44557 37247
rect 42852 37216 44557 37244
rect 42852 37204 42858 37216
rect 44545 37213 44557 37216
rect 44591 37213 44603 37247
rect 44545 37207 44603 37213
rect 45465 37247 45523 37253
rect 45465 37213 45477 37247
rect 45511 37244 45523 37247
rect 45738 37244 45744 37256
rect 45511 37216 45744 37244
rect 45511 37213 45523 37216
rect 45465 37207 45523 37213
rect 45738 37204 45744 37216
rect 45796 37204 45802 37256
rect 47210 37204 47216 37256
rect 47268 37204 47274 37256
rect 47504 37244 47532 37284
rect 49789 37281 49801 37284
rect 49835 37312 49847 37315
rect 50341 37315 50399 37321
rect 50341 37312 50353 37315
rect 49835 37284 50353 37312
rect 49835 37281 49847 37284
rect 49789 37275 49847 37281
rect 50341 37281 50353 37284
rect 50387 37281 50399 37315
rect 52914 37312 52920 37324
rect 50341 37275 50399 37281
rect 52472 37284 52920 37312
rect 47320 37216 47532 37244
rect 47949 37247 48007 37253
rect 30340 37148 31754 37176
rect 30340 37136 30346 37148
rect 46750 37136 46756 37188
rect 46808 37176 46814 37188
rect 47320 37176 47348 37216
rect 47949 37213 47961 37247
rect 47995 37213 48007 37247
rect 47949 37207 48007 37213
rect 48133 37247 48191 37253
rect 48133 37213 48145 37247
rect 48179 37244 48191 37247
rect 48179 37216 48314 37244
rect 48179 37213 48191 37216
rect 48133 37207 48191 37213
rect 46808 37148 47348 37176
rect 46808 37136 46814 37148
rect 18555 37080 18828 37108
rect 18555 37077 18567 37080
rect 18509 37071 18567 37077
rect 26970 37068 26976 37120
rect 27028 37108 27034 37120
rect 38654 37108 38660 37120
rect 27028 37080 38660 37108
rect 27028 37068 27034 37080
rect 38654 37068 38660 37080
rect 38712 37068 38718 37120
rect 41690 37068 41696 37120
rect 41748 37068 41754 37120
rect 47118 37068 47124 37120
rect 47176 37108 47182 37120
rect 47964 37108 47992 37207
rect 48286 37176 48314 37216
rect 48590 37204 48596 37256
rect 48648 37244 48654 37256
rect 50525 37247 50583 37253
rect 50525 37244 50537 37247
rect 48648 37216 50537 37244
rect 48648 37204 48654 37216
rect 50525 37213 50537 37216
rect 50571 37213 50583 37247
rect 50525 37207 50583 37213
rect 51537 37247 51595 37253
rect 51537 37213 51549 37247
rect 51583 37244 51595 37247
rect 52472 37244 52500 37284
rect 52914 37272 52920 37284
rect 52972 37272 52978 37324
rect 53576 37284 53788 37312
rect 53576 37253 53604 37284
rect 51583 37216 52500 37244
rect 52825 37247 52883 37253
rect 51583 37213 51595 37216
rect 51537 37207 51595 37213
rect 52825 37213 52837 37247
rect 52871 37213 52883 37247
rect 52825 37207 52883 37213
rect 53561 37247 53619 37253
rect 53561 37213 53573 37247
rect 53607 37213 53619 37247
rect 53561 37207 53619 37213
rect 53653 37247 53711 37253
rect 53653 37213 53665 37247
rect 53699 37213 53711 37247
rect 53760 37244 53788 37284
rect 56042 37272 56048 37324
rect 56100 37272 56106 37324
rect 57146 37272 57152 37324
rect 57204 37312 57210 37324
rect 57609 37315 57667 37321
rect 57609 37312 57621 37315
rect 57204 37284 57621 37312
rect 57204 37272 57210 37284
rect 57609 37281 57621 37284
rect 57655 37281 57667 37315
rect 57609 37275 57667 37281
rect 58986 37272 58992 37324
rect 59044 37272 59050 37324
rect 59188 37312 59216 37420
rect 59262 37408 59268 37460
rect 59320 37448 59326 37460
rect 59320 37420 60734 37448
rect 59320 37408 59326 37420
rect 59633 37383 59691 37389
rect 59633 37349 59645 37383
rect 59679 37380 59691 37383
rect 59814 37380 59820 37392
rect 59679 37352 59820 37380
rect 59679 37349 59691 37352
rect 59633 37343 59691 37349
rect 59814 37340 59820 37352
rect 59872 37340 59878 37392
rect 60706 37380 60734 37420
rect 62482 37408 62488 37460
rect 62540 37408 62546 37460
rect 65794 37448 65800 37460
rect 62684 37420 65800 37448
rect 62684 37380 62712 37420
rect 65794 37408 65800 37420
rect 65852 37408 65858 37460
rect 60706 37352 62790 37380
rect 62482 37312 62488 37324
rect 59188 37284 62488 37312
rect 62482 37272 62488 37284
rect 62540 37272 62546 37324
rect 64230 37272 64236 37324
rect 64288 37272 64294 37324
rect 56226 37244 56232 37256
rect 53760 37216 56232 37244
rect 53653 37207 53711 37213
rect 48682 37176 48688 37188
rect 48286 37148 48688 37176
rect 48682 37136 48688 37148
rect 48740 37136 48746 37188
rect 47176 37080 47992 37108
rect 52840 37108 52868 37207
rect 53190 37136 53196 37188
rect 53248 37176 53254 37188
rect 53668 37176 53696 37207
rect 56226 37204 56232 37216
rect 56284 37204 56290 37256
rect 56594 37204 56600 37256
rect 56652 37204 56658 37256
rect 57885 37247 57943 37253
rect 57885 37244 57897 37247
rect 57164 37216 57897 37244
rect 53742 37176 53748 37188
rect 53248 37148 53748 37176
rect 53248 37136 53254 37148
rect 53742 37136 53748 37148
rect 53800 37136 53806 37188
rect 57164 37185 57192 37216
rect 57885 37213 57897 37216
rect 57931 37213 57943 37247
rect 57885 37207 57943 37213
rect 63862 37204 63868 37256
rect 63920 37244 63926 37256
rect 63957 37247 64015 37253
rect 63957 37244 63969 37247
rect 63920 37216 63969 37244
rect 63920 37204 63926 37216
rect 63957 37213 63969 37216
rect 64003 37213 64015 37247
rect 63957 37207 64015 37213
rect 65702 37204 65708 37256
rect 65760 37244 65766 37256
rect 65981 37247 66039 37253
rect 65981 37244 65993 37247
rect 65760 37216 65993 37244
rect 65760 37204 65766 37216
rect 65981 37213 65993 37216
rect 66027 37213 66039 37247
rect 65981 37207 66039 37213
rect 57149 37179 57207 37185
rect 57149 37145 57161 37179
rect 57195 37145 57207 37179
rect 57149 37139 57207 37145
rect 54662 37108 54668 37120
rect 52840 37080 54668 37108
rect 47176 37068 47182 37080
rect 54662 37068 54668 37080
rect 54720 37068 54726 37120
rect 65426 37068 65432 37120
rect 65484 37068 65490 37120
rect 552 37018 66424 37040
rect 552 36966 1998 37018
rect 2050 36966 2062 37018
rect 2114 36966 2126 37018
rect 2178 36966 2190 37018
rect 2242 36966 2254 37018
rect 2306 36966 49998 37018
rect 50050 36966 50062 37018
rect 50114 36966 50126 37018
rect 50178 36966 50190 37018
rect 50242 36966 50254 37018
rect 50306 36966 64338 37018
rect 64390 36966 64402 37018
rect 64454 36966 64466 37018
rect 64518 36966 64530 37018
rect 64582 36966 64594 37018
rect 64646 36966 66424 37018
rect 552 36944 66424 36966
rect 23474 36864 23480 36916
rect 23532 36904 23538 36916
rect 28994 36904 29000 36916
rect 23532 36876 29000 36904
rect 23532 36864 23538 36876
rect 28994 36864 29000 36876
rect 29052 36864 29058 36916
rect 31294 36864 31300 36916
rect 31352 36904 31358 36916
rect 35710 36904 35716 36916
rect 31352 36876 35716 36904
rect 31352 36864 31358 36876
rect 35710 36864 35716 36876
rect 35768 36864 35774 36916
rect 42242 36864 42248 36916
rect 42300 36904 42306 36916
rect 42300 36876 44220 36904
rect 42300 36864 42306 36876
rect 21174 36796 21180 36848
rect 21232 36836 21238 36848
rect 44082 36836 44088 36848
rect 21232 36808 44088 36836
rect 21232 36796 21238 36808
rect 44082 36796 44088 36808
rect 44140 36796 44146 36848
rect 44192 36836 44220 36876
rect 47210 36864 47216 36916
rect 47268 36904 47274 36916
rect 48590 36904 48596 36916
rect 47268 36876 48596 36904
rect 47268 36864 47274 36876
rect 48590 36864 48596 36876
rect 48648 36864 48654 36916
rect 62850 36904 62856 36916
rect 51046 36876 62856 36904
rect 51046 36836 51074 36876
rect 62850 36864 62856 36876
rect 62908 36864 62914 36916
rect 63862 36864 63868 36916
rect 63920 36864 63926 36916
rect 66162 36836 66168 36848
rect 44192 36808 51074 36836
rect 57946 36808 66168 36836
rect 22002 36728 22008 36780
rect 22060 36768 22066 36780
rect 46750 36768 46756 36780
rect 22060 36740 46756 36768
rect 22060 36728 22066 36740
rect 46750 36728 46756 36740
rect 46808 36728 46814 36780
rect 38838 36660 38844 36712
rect 38896 36700 38902 36712
rect 57946 36700 57974 36808
rect 66162 36796 66168 36808
rect 66220 36796 66226 36848
rect 60642 36728 60648 36780
rect 60700 36768 60706 36780
rect 64417 36771 64475 36777
rect 64417 36768 64429 36771
rect 60700 36740 64429 36768
rect 60700 36728 60706 36740
rect 64417 36737 64429 36740
rect 64463 36768 64475 36771
rect 65245 36771 65303 36777
rect 65245 36768 65257 36771
rect 64463 36740 65257 36768
rect 64463 36737 64475 36740
rect 64417 36731 64475 36737
rect 65245 36737 65257 36740
rect 65291 36768 65303 36771
rect 66530 36768 66536 36780
rect 65291 36740 66536 36768
rect 65291 36737 65303 36740
rect 65245 36731 65303 36737
rect 66530 36728 66536 36740
rect 66588 36728 66594 36780
rect 38896 36672 57974 36700
rect 38896 36660 38902 36672
rect 64046 36660 64052 36712
rect 64104 36700 64110 36712
rect 64233 36703 64291 36709
rect 64233 36700 64245 36703
rect 64104 36672 64245 36700
rect 64104 36660 64110 36672
rect 64233 36669 64245 36672
rect 64279 36669 64291 36703
rect 64233 36663 64291 36669
rect 65061 36703 65119 36709
rect 65061 36669 65073 36703
rect 65107 36700 65119 36703
rect 65426 36700 65432 36712
rect 65107 36672 65432 36700
rect 65107 36669 65119 36672
rect 65061 36663 65119 36669
rect 65426 36660 65432 36672
rect 65484 36660 65490 36712
rect 24854 36592 24860 36644
rect 24912 36632 24918 36644
rect 34422 36632 34428 36644
rect 24912 36604 34428 36632
rect 24912 36592 24918 36604
rect 34422 36592 34428 36604
rect 34480 36592 34486 36644
rect 37274 36592 37280 36644
rect 37332 36632 37338 36644
rect 64325 36635 64383 36641
rect 37332 36604 55996 36632
rect 37332 36592 37338 36604
rect 11698 36524 11704 36576
rect 11756 36564 11762 36576
rect 11756 36536 55904 36564
rect 11756 36524 11762 36536
rect 8478 36456 8484 36508
rect 8536 36496 8542 36508
rect 52546 36496 52552 36508
rect 8536 36468 52552 36496
rect 8536 36456 8542 36468
rect 52546 36456 52552 36468
rect 52604 36456 52610 36508
rect 21542 36388 21548 36440
rect 21600 36428 21606 36440
rect 28994 36428 29000 36440
rect 21600 36400 29000 36428
rect 21600 36388 21606 36400
rect 28994 36388 29000 36400
rect 29052 36388 29058 36440
rect 30282 36320 30288 36372
rect 30340 36360 30346 36372
rect 33042 36360 33048 36372
rect 30340 36332 33048 36360
rect 30340 36320 30346 36332
rect 33042 36320 33048 36332
rect 33100 36320 33106 36372
rect 44082 36252 44088 36304
rect 44140 36292 44146 36304
rect 55876 36292 55904 36536
rect 55968 36360 55996 36604
rect 64325 36601 64337 36635
rect 64371 36632 64383 36635
rect 64782 36632 64788 36644
rect 64371 36604 64788 36632
rect 64371 36601 64383 36604
rect 64325 36595 64383 36601
rect 64782 36592 64788 36604
rect 64840 36592 64846 36644
rect 64138 36524 64144 36576
rect 64196 36564 64202 36576
rect 64693 36567 64751 36573
rect 64693 36564 64705 36567
rect 64196 36536 64705 36564
rect 64196 36524 64202 36536
rect 64693 36533 64705 36536
rect 64739 36533 64751 36567
rect 64693 36527 64751 36533
rect 65150 36524 65156 36576
rect 65208 36524 65214 36576
rect 63572 36474 66424 36496
rect 63572 36422 65258 36474
rect 65310 36422 65322 36474
rect 65374 36422 65386 36474
rect 65438 36422 65450 36474
rect 65502 36422 65514 36474
rect 65566 36422 66424 36474
rect 63572 36400 66424 36422
rect 66070 36360 66076 36372
rect 55968 36332 66076 36360
rect 66070 36320 66076 36332
rect 66128 36320 66134 36372
rect 61562 36292 61568 36304
rect 44140 36264 51074 36292
rect 55876 36264 61568 36292
rect 44140 36252 44146 36264
rect 25866 36184 25872 36236
rect 25924 36224 25930 36236
rect 51046 36224 51074 36264
rect 61562 36252 61568 36264
rect 61620 36252 61626 36304
rect 63218 36252 63224 36304
rect 63276 36292 63282 36304
rect 63494 36292 63500 36304
rect 63276 36264 63500 36292
rect 63276 36252 63282 36264
rect 63494 36252 63500 36264
rect 63552 36252 63558 36304
rect 64138 36252 64144 36304
rect 64196 36252 64202 36304
rect 65794 36292 65800 36304
rect 65366 36264 65800 36292
rect 65794 36252 65800 36264
rect 65852 36252 65858 36304
rect 63678 36224 63684 36236
rect 25924 36196 44680 36224
rect 51046 36196 63684 36224
rect 25924 36184 25930 36196
rect 27614 36116 27620 36168
rect 27672 36156 27678 36168
rect 43530 36156 43536 36168
rect 27672 36128 43536 36156
rect 27672 36116 27678 36128
rect 43530 36116 43536 36128
rect 43588 36116 43594 36168
rect 44652 36156 44680 36196
rect 63678 36184 63684 36196
rect 63736 36184 63742 36236
rect 63770 36156 63776 36168
rect 44652 36128 63776 36156
rect 63770 36116 63776 36128
rect 63828 36116 63834 36168
rect 63862 36116 63868 36168
rect 63920 36116 63926 36168
rect 23198 36048 23204 36100
rect 23256 36088 23262 36100
rect 38654 36088 38660 36100
rect 23256 36060 38660 36088
rect 23256 36048 23262 36060
rect 38654 36048 38660 36060
rect 38712 36048 38718 36100
rect 24670 35980 24676 36032
rect 24728 36020 24734 36032
rect 28534 36020 28540 36032
rect 24728 35992 28540 36020
rect 24728 35980 24734 35992
rect 28534 35980 28540 35992
rect 28592 35980 28598 36032
rect 29086 35980 29092 36032
rect 29144 36020 29150 36032
rect 62574 36020 62580 36032
rect 29144 35992 62580 36020
rect 29144 35980 29150 35992
rect 62574 35980 62580 35992
rect 62632 35980 62638 36032
rect 65613 36023 65671 36029
rect 65613 35989 65625 36023
rect 65659 36020 65671 36023
rect 65702 36020 65708 36032
rect 65659 35992 65708 36020
rect 65659 35989 65671 35992
rect 65613 35983 65671 35989
rect 65702 35980 65708 35992
rect 65760 35980 65766 36032
rect 35802 35952 35808 35964
rect 29012 35924 35808 35952
rect 20070 35844 20076 35896
rect 20128 35884 20134 35896
rect 23106 35884 23112 35896
rect 20128 35856 23112 35884
rect 20128 35844 20134 35856
rect 23106 35844 23112 35856
rect 23164 35844 23170 35896
rect 23566 35844 23572 35896
rect 23624 35884 23630 35896
rect 29012 35884 29040 35924
rect 35802 35912 35808 35924
rect 35860 35912 35866 35964
rect 63572 35930 66424 35952
rect 23624 35856 29040 35884
rect 23624 35844 23630 35856
rect 30006 35844 30012 35896
rect 30064 35884 30070 35896
rect 44082 35884 44088 35896
rect 30064 35856 44088 35884
rect 30064 35844 30070 35856
rect 44082 35844 44088 35856
rect 44140 35844 44146 35896
rect 63572 35878 64338 35930
rect 64390 35878 64402 35930
rect 64454 35878 64466 35930
rect 64518 35878 64530 35930
rect 64582 35878 64594 35930
rect 64646 35878 66424 35930
rect 63572 35856 66424 35878
rect 28994 35776 29000 35828
rect 29052 35816 29058 35828
rect 33134 35816 33140 35828
rect 29052 35788 33140 35816
rect 29052 35776 29058 35788
rect 33134 35776 33140 35788
rect 33192 35776 33198 35828
rect 35710 35776 35716 35828
rect 35768 35816 35774 35828
rect 40034 35816 40040 35828
rect 35768 35788 40040 35816
rect 35768 35776 35774 35788
rect 40034 35776 40040 35788
rect 40092 35776 40098 35828
rect 60550 35776 60556 35828
rect 60608 35816 60614 35828
rect 65061 35819 65119 35825
rect 60608 35788 63816 35816
rect 60608 35776 60614 35788
rect 23014 35708 23020 35760
rect 23072 35748 23078 35760
rect 29086 35748 29092 35760
rect 23072 35720 29092 35748
rect 23072 35708 23078 35720
rect 29086 35708 29092 35720
rect 29144 35708 29150 35760
rect 31570 35708 31576 35760
rect 31628 35748 31634 35760
rect 33594 35748 33600 35760
rect 31628 35720 33600 35748
rect 31628 35708 31634 35720
rect 33594 35708 33600 35720
rect 33652 35708 33658 35760
rect 63586 35640 63592 35692
rect 63644 35640 63650 35692
rect 63788 35680 63816 35788
rect 65061 35785 65073 35819
rect 65107 35816 65119 35819
rect 65150 35816 65156 35828
rect 65107 35788 65156 35816
rect 65107 35785 65119 35788
rect 65061 35779 65119 35785
rect 65150 35776 65156 35788
rect 65208 35776 65214 35828
rect 63954 35708 63960 35760
rect 64012 35748 64018 35760
rect 64012 35720 65196 35748
rect 64012 35708 64018 35720
rect 65168 35692 65196 35720
rect 64785 35683 64843 35689
rect 64785 35680 64797 35683
rect 63788 35652 64797 35680
rect 64785 35649 64797 35652
rect 64831 35649 64843 35683
rect 64785 35643 64843 35649
rect 65150 35640 65156 35692
rect 65208 35640 65214 35692
rect 65518 35640 65524 35692
rect 65576 35640 65582 35692
rect 65610 35640 65616 35692
rect 65668 35640 65674 35692
rect 61562 35572 61568 35624
rect 61620 35612 61626 35624
rect 62482 35612 62488 35624
rect 61620 35584 62488 35612
rect 61620 35572 61626 35584
rect 62482 35572 62488 35584
rect 62540 35572 62546 35624
rect 63604 35612 63632 35640
rect 63770 35612 63776 35624
rect 63604 35584 63776 35612
rect 63770 35572 63776 35584
rect 63828 35572 63834 35624
rect 63954 35572 63960 35624
rect 64012 35612 64018 35624
rect 64601 35615 64659 35621
rect 64601 35612 64613 35615
rect 64012 35584 64613 35612
rect 64012 35572 64018 35584
rect 64601 35581 64613 35584
rect 64647 35581 64659 35615
rect 64601 35575 64659 35581
rect 8202 35504 8208 35556
rect 8260 35544 8266 35556
rect 18046 35544 18052 35556
rect 8260 35516 18052 35544
rect 8260 35504 8266 35516
rect 18046 35504 18052 35516
rect 18104 35504 18110 35556
rect 22186 35504 22192 35556
rect 22244 35544 22250 35556
rect 64046 35544 64052 35556
rect 22244 35516 64052 35544
rect 22244 35504 22250 35516
rect 64046 35504 64052 35516
rect 64104 35504 64110 35556
rect 65429 35547 65487 35553
rect 65429 35513 65441 35547
rect 65475 35544 65487 35547
rect 65978 35544 65984 35556
rect 65475 35516 65984 35544
rect 65475 35513 65487 35516
rect 65429 35507 65487 35513
rect 65978 35504 65984 35516
rect 66036 35504 66042 35556
rect 64138 35436 64144 35488
rect 64196 35476 64202 35488
rect 64233 35479 64291 35485
rect 64233 35476 64245 35479
rect 64196 35448 64245 35476
rect 64196 35436 64202 35448
rect 64233 35445 64245 35448
rect 64279 35445 64291 35479
rect 64233 35439 64291 35445
rect 64690 35436 64696 35488
rect 64748 35436 64754 35488
rect 63572 35386 66424 35408
rect 63572 35334 65258 35386
rect 65310 35334 65322 35386
rect 65374 35334 65386 35386
rect 65438 35334 65450 35386
rect 65502 35334 65514 35386
rect 65566 35334 66424 35386
rect 63572 35312 66424 35334
rect 62942 35232 62948 35284
rect 63000 35272 63006 35284
rect 65610 35272 65616 35284
rect 63000 35244 65616 35272
rect 63000 35232 63006 35244
rect 65610 35232 65616 35244
rect 65668 35272 65674 35284
rect 65886 35272 65892 35284
rect 65668 35244 65892 35272
rect 65668 35232 65674 35244
rect 65886 35232 65892 35244
rect 65944 35232 65950 35284
rect 64138 35164 64144 35216
rect 64196 35164 64202 35216
rect 65794 35204 65800 35216
rect 65366 35176 65800 35204
rect 65794 35164 65800 35176
rect 65852 35164 65858 35216
rect 63862 35028 63868 35080
rect 63920 35028 63926 35080
rect 64138 35028 64144 35080
rect 64196 35068 64202 35080
rect 64598 35068 64604 35080
rect 64196 35040 64604 35068
rect 64196 35028 64202 35040
rect 64598 35028 64604 35040
rect 64656 35028 64662 35080
rect 63880 34932 63908 35028
rect 65150 34932 65156 34944
rect 63880 34904 65156 34932
rect 65150 34892 65156 34904
rect 65208 34892 65214 34944
rect 65610 34892 65616 34944
rect 65668 34892 65674 34944
rect 63572 34842 66424 34864
rect 63572 34790 64338 34842
rect 64390 34790 64402 34842
rect 64454 34790 64466 34842
rect 64518 34790 64530 34842
rect 64582 34790 64594 34842
rect 64646 34790 66424 34842
rect 63572 34768 66424 34790
rect 64690 34688 64696 34740
rect 64748 34688 64754 34740
rect 64601 34663 64659 34669
rect 64156 34632 64552 34660
rect 62942 34552 62948 34604
rect 63000 34592 63006 34604
rect 63957 34595 64015 34601
rect 63957 34592 63969 34595
rect 63000 34564 63969 34592
rect 63000 34552 63006 34564
rect 63957 34561 63969 34564
rect 64003 34561 64015 34595
rect 63957 34555 64015 34561
rect 64156 34533 64184 34632
rect 64141 34527 64199 34533
rect 64141 34493 64153 34527
rect 64187 34493 64199 34527
rect 64524 34524 64552 34632
rect 64601 34629 64613 34663
rect 64647 34660 64659 34663
rect 64782 34660 64788 34672
rect 64647 34632 64788 34660
rect 64647 34629 64659 34632
rect 64601 34623 64659 34629
rect 64782 34620 64788 34632
rect 64840 34620 64846 34672
rect 66254 34660 66260 34672
rect 65168 34632 66260 34660
rect 65168 34601 65196 34632
rect 66254 34620 66260 34632
rect 66312 34620 66318 34672
rect 65153 34595 65211 34601
rect 65153 34561 65165 34595
rect 65199 34561 65211 34595
rect 65153 34555 65211 34561
rect 65242 34552 65248 34604
rect 65300 34552 65306 34604
rect 65610 34524 65616 34536
rect 64524 34496 65616 34524
rect 64141 34487 64199 34493
rect 65610 34484 65616 34496
rect 65668 34484 65674 34536
rect 64046 34416 64052 34468
rect 64104 34456 64110 34468
rect 64233 34459 64291 34465
rect 64233 34456 64245 34459
rect 64104 34428 64245 34456
rect 64104 34416 64110 34428
rect 64233 34425 64245 34428
rect 64279 34425 64291 34459
rect 64233 34419 64291 34425
rect 64322 34416 64328 34468
rect 64380 34456 64386 34468
rect 65061 34459 65119 34465
rect 65061 34456 65073 34459
rect 64380 34428 65073 34456
rect 64380 34416 64386 34428
rect 65061 34425 65073 34428
rect 65107 34425 65119 34459
rect 65061 34419 65119 34425
rect 63678 34348 63684 34400
rect 63736 34388 63742 34400
rect 64782 34388 64788 34400
rect 63736 34360 64788 34388
rect 63736 34348 63742 34360
rect 64782 34348 64788 34360
rect 64840 34348 64846 34400
rect 63572 34298 66424 34320
rect 63572 34246 65258 34298
rect 65310 34246 65322 34298
rect 65374 34246 65386 34298
rect 65438 34246 65450 34298
rect 65502 34246 65514 34298
rect 65566 34246 66424 34298
rect 63572 34224 66424 34246
rect 63954 34144 63960 34196
rect 64012 34184 64018 34196
rect 65153 34187 65211 34193
rect 65153 34184 65165 34187
rect 64012 34156 65165 34184
rect 64012 34144 64018 34156
rect 65153 34153 65165 34156
rect 65199 34153 65211 34187
rect 65153 34147 65211 34153
rect 63402 34076 63408 34128
rect 63460 34116 63466 34128
rect 64322 34116 64328 34128
rect 63460 34088 64328 34116
rect 63460 34076 63466 34088
rect 64322 34076 64328 34088
rect 64380 34076 64386 34128
rect 65610 34008 65616 34060
rect 65668 34048 65674 34060
rect 65705 34051 65763 34057
rect 65705 34048 65717 34051
rect 65668 34020 65717 34048
rect 65668 34008 65674 34020
rect 65705 34017 65717 34020
rect 65751 34017 65763 34051
rect 65705 34011 65763 34017
rect 63218 33940 63224 33992
rect 63276 33980 63282 33992
rect 64138 33980 64144 33992
rect 63276 33952 64144 33980
rect 63276 33940 63282 33952
rect 64138 33940 64144 33952
rect 64196 33940 64202 33992
rect 63770 33804 63776 33856
rect 63828 33844 63834 33856
rect 64966 33844 64972 33856
rect 63828 33816 64972 33844
rect 63828 33804 63834 33816
rect 64966 33804 64972 33816
rect 65024 33804 65030 33856
rect 63572 33754 66424 33776
rect 63572 33702 64338 33754
rect 64390 33702 64402 33754
rect 64454 33702 64466 33754
rect 64518 33702 64530 33754
rect 64582 33702 64594 33754
rect 64646 33702 66424 33754
rect 63572 33680 66424 33702
rect 66530 33572 66536 33584
rect 65168 33544 66536 33572
rect 65168 33513 65196 33544
rect 66530 33532 66536 33544
rect 66588 33532 66594 33584
rect 65153 33507 65211 33513
rect 65153 33473 65165 33507
rect 65199 33473 65211 33507
rect 65153 33467 65211 33473
rect 65978 33464 65984 33516
rect 66036 33464 66042 33516
rect 64877 33371 64935 33377
rect 64877 33337 64889 33371
rect 64923 33368 64935 33371
rect 65429 33371 65487 33377
rect 65429 33368 65441 33371
rect 64923 33340 65441 33368
rect 64923 33337 64935 33340
rect 64877 33331 64935 33337
rect 65429 33337 65441 33340
rect 65475 33337 65487 33371
rect 65429 33331 65487 33337
rect 64322 33260 64328 33312
rect 64380 33300 64386 33312
rect 64509 33303 64567 33309
rect 64509 33300 64521 33303
rect 64380 33272 64521 33300
rect 64380 33260 64386 33272
rect 64509 33269 64521 33272
rect 64555 33269 64567 33303
rect 64509 33263 64567 33269
rect 64966 33260 64972 33312
rect 65024 33260 65030 33312
rect 63572 33210 66424 33232
rect 63572 33158 65258 33210
rect 65310 33158 65322 33210
rect 65374 33158 65386 33210
rect 65438 33158 65450 33210
rect 65502 33158 65514 33210
rect 65566 33158 66424 33210
rect 63572 33136 66424 33158
rect 65797 33099 65855 33105
rect 65797 33065 65809 33099
rect 65843 33096 65855 33099
rect 65978 33096 65984 33108
rect 65843 33068 65984 33096
rect 65843 33065 65855 33068
rect 65797 33059 65855 33065
rect 65978 33056 65984 33068
rect 66036 33056 66042 33108
rect 64230 33028 64236 33040
rect 64064 33000 64236 33028
rect 64064 32972 64092 33000
rect 64230 32988 64236 33000
rect 64288 32988 64294 33040
rect 64322 32988 64328 33040
rect 64380 32988 64386 33040
rect 66346 33028 66352 33040
rect 65550 33000 66352 33028
rect 66346 32988 66352 33000
rect 66404 32988 66410 33040
rect 64046 32920 64052 32972
rect 64104 32920 64110 32972
rect 63572 32666 66424 32688
rect 63572 32614 64338 32666
rect 64390 32614 64402 32666
rect 64454 32614 64466 32666
rect 64518 32614 64530 32666
rect 64582 32614 64594 32666
rect 64646 32614 66424 32666
rect 63572 32592 66424 32614
rect 64966 32512 64972 32564
rect 65024 32552 65030 32564
rect 65061 32555 65119 32561
rect 65061 32552 65073 32555
rect 65024 32524 65073 32552
rect 65024 32512 65030 32524
rect 65061 32521 65073 32524
rect 65107 32521 65119 32555
rect 65061 32515 65119 32521
rect 65886 32484 65892 32496
rect 64524 32456 65892 32484
rect 64524 32425 64552 32456
rect 65886 32444 65892 32456
rect 65944 32444 65950 32496
rect 64509 32419 64567 32425
rect 64509 32385 64521 32419
rect 64555 32385 64567 32419
rect 64509 32379 64567 32385
rect 64601 32419 64659 32425
rect 64601 32385 64613 32419
rect 64647 32416 64659 32419
rect 65702 32416 65708 32428
rect 64647 32388 65708 32416
rect 64647 32385 64659 32388
rect 64601 32379 64659 32385
rect 65702 32376 65708 32388
rect 65760 32376 65766 32428
rect 64690 32308 64696 32360
rect 64748 32308 64754 32360
rect 64966 32172 64972 32224
rect 65024 32212 65030 32224
rect 65978 32212 65984 32224
rect 65024 32184 65984 32212
rect 65024 32172 65030 32184
rect 65978 32172 65984 32184
rect 66036 32172 66042 32224
rect 63572 32122 66424 32144
rect 63572 32070 65258 32122
rect 65310 32070 65322 32122
rect 65374 32070 65386 32122
rect 65438 32070 65450 32122
rect 65502 32070 65514 32122
rect 65566 32070 66424 32122
rect 63572 32048 66424 32070
rect 64969 32011 65027 32017
rect 64969 31977 64981 32011
rect 65015 32008 65027 32011
rect 65337 32011 65395 32017
rect 65015 31980 65288 32008
rect 65015 31977 65027 31980
rect 64969 31971 65027 31977
rect 65260 31940 65288 31980
rect 65337 31977 65349 32011
rect 65383 32008 65395 32011
rect 65794 32008 65800 32020
rect 65383 31980 65800 32008
rect 65383 31977 65395 31980
rect 65337 31971 65395 31977
rect 65794 31968 65800 31980
rect 65852 31968 65858 32020
rect 65610 31940 65616 31952
rect 64800 31912 65104 31940
rect 65260 31912 65616 31940
rect 64800 31813 64828 31912
rect 64877 31875 64935 31881
rect 64877 31841 64889 31875
rect 64923 31872 64935 31875
rect 64966 31872 64972 31884
rect 64923 31844 64972 31872
rect 64923 31841 64935 31844
rect 64877 31835 64935 31841
rect 64966 31832 64972 31844
rect 65024 31832 65030 31884
rect 64785 31807 64843 31813
rect 64785 31773 64797 31807
rect 64831 31773 64843 31807
rect 65076 31804 65104 31912
rect 65610 31900 65616 31912
rect 65668 31900 65674 31952
rect 65334 31832 65340 31884
rect 65392 31872 65398 31884
rect 65886 31872 65892 31884
rect 65392 31844 65892 31872
rect 65392 31832 65398 31844
rect 65886 31832 65892 31844
rect 65944 31832 65950 31884
rect 66438 31832 66444 31884
rect 66496 31832 66502 31884
rect 65242 31804 65248 31816
rect 64785 31767 64843 31773
rect 64984 31776 65248 31804
rect 64984 31748 65012 31776
rect 65242 31764 65248 31776
rect 65300 31764 65306 31816
rect 65521 31807 65579 31813
rect 65521 31773 65533 31807
rect 65567 31804 65579 31807
rect 65567 31776 65656 31804
rect 65567 31773 65579 31776
rect 65521 31767 65579 31773
rect 64966 31696 64972 31748
rect 65024 31696 65030 31748
rect 65628 31736 65656 31776
rect 65702 31764 65708 31816
rect 65760 31804 65766 31816
rect 66073 31807 66131 31813
rect 66073 31804 66085 31807
rect 65760 31776 66085 31804
rect 65760 31764 65766 31776
rect 66073 31773 66085 31776
rect 66119 31773 66131 31807
rect 66073 31767 66131 31773
rect 66162 31764 66168 31816
rect 66220 31804 66226 31816
rect 66456 31804 66484 31832
rect 66220 31776 66484 31804
rect 66220 31764 66226 31776
rect 65978 31736 65984 31748
rect 65628 31708 65984 31736
rect 65978 31696 65984 31708
rect 66036 31696 66042 31748
rect 63572 31578 66424 31600
rect 63572 31526 64338 31578
rect 64390 31526 64402 31578
rect 64454 31526 64466 31578
rect 64518 31526 64530 31578
rect 64582 31526 64594 31578
rect 64646 31526 66424 31578
rect 63572 31504 66424 31526
rect 64046 31424 64052 31476
rect 64104 31464 64110 31476
rect 65153 31467 65211 31473
rect 65153 31464 65165 31467
rect 64104 31436 65165 31464
rect 64104 31424 64110 31436
rect 65153 31433 65165 31436
rect 65199 31433 65211 31467
rect 65153 31427 65211 31433
rect 63865 31263 63923 31269
rect 63865 31229 63877 31263
rect 63911 31260 63923 31263
rect 64966 31260 64972 31272
rect 63911 31232 64972 31260
rect 63911 31229 63923 31232
rect 63865 31223 63923 31229
rect 64966 31220 64972 31232
rect 65024 31220 65030 31272
rect 65058 31220 65064 31272
rect 65116 31260 65122 31272
rect 65242 31260 65248 31272
rect 65116 31232 65248 31260
rect 65116 31220 65122 31232
rect 65242 31220 65248 31232
rect 65300 31220 65306 31272
rect 63572 31034 66424 31056
rect 63572 30982 65258 31034
rect 65310 30982 65322 31034
rect 65374 30982 65386 31034
rect 65438 30982 65450 31034
rect 65502 30982 65514 31034
rect 65566 30982 66424 31034
rect 63572 30960 66424 30982
rect 65150 30880 65156 30932
rect 65208 30880 65214 30932
rect 63862 30744 63868 30796
rect 63920 30784 63926 30796
rect 64874 30784 64880 30796
rect 63920 30756 64880 30784
rect 63920 30744 63926 30756
rect 64874 30744 64880 30756
rect 64932 30744 64938 30796
rect 64874 30608 64880 30660
rect 64932 30648 64938 30660
rect 65058 30648 65064 30660
rect 64932 30620 65064 30648
rect 64932 30608 64938 30620
rect 65058 30608 65064 30620
rect 65116 30608 65122 30660
rect 63572 30490 66424 30512
rect 63572 30438 64338 30490
rect 64390 30438 64402 30490
rect 64454 30438 64466 30490
rect 64518 30438 64530 30490
rect 64582 30438 64594 30490
rect 64646 30438 66424 30490
rect 63572 30416 66424 30438
rect 64049 30243 64107 30249
rect 64049 30209 64061 30243
rect 64095 30240 64107 30243
rect 65058 30240 65064 30252
rect 64095 30212 65064 30240
rect 64095 30209 64107 30212
rect 64049 30203 64107 30209
rect 65058 30200 65064 30212
rect 65116 30200 65122 30252
rect 64322 30064 64328 30116
rect 64380 30064 64386 30116
rect 66438 30104 66444 30116
rect 65550 30076 66444 30104
rect 66438 30064 66444 30076
rect 66496 30064 66502 30116
rect 65797 30039 65855 30045
rect 65797 30005 65809 30039
rect 65843 30036 65855 30039
rect 65978 30036 65984 30048
rect 65843 30008 65984 30036
rect 65843 30005 65855 30008
rect 65797 29999 65855 30005
rect 65978 29996 65984 30008
rect 66036 29996 66042 30048
rect 62942 29928 62948 29980
rect 63000 29968 63006 29980
rect 63126 29968 63132 29980
rect 63000 29940 63132 29968
rect 63000 29928 63006 29940
rect 63126 29928 63132 29940
rect 63184 29928 63190 29980
rect 63572 29946 66424 29968
rect 63572 29894 65258 29946
rect 65310 29894 65322 29946
rect 65374 29894 65386 29946
rect 65438 29894 65450 29946
rect 65502 29894 65514 29946
rect 65566 29894 66424 29946
rect 63572 29872 66424 29894
rect 64322 29792 64328 29844
rect 64380 29832 64386 29844
rect 65337 29835 65395 29841
rect 65337 29832 65349 29835
rect 64380 29804 65349 29832
rect 64380 29792 64386 29804
rect 65337 29801 65349 29804
rect 65383 29801 65395 29835
rect 65337 29795 65395 29801
rect 65702 29792 65708 29844
rect 65760 29792 65766 29844
rect 65794 29792 65800 29844
rect 65852 29792 65858 29844
rect 64877 29767 64935 29773
rect 64877 29733 64889 29767
rect 64923 29764 64935 29767
rect 65058 29764 65064 29776
rect 64923 29736 65064 29764
rect 64923 29733 64935 29736
rect 64877 29727 64935 29733
rect 65058 29724 65064 29736
rect 65116 29724 65122 29776
rect 64969 29699 65027 29705
rect 64969 29665 64981 29699
rect 65015 29696 65027 29699
rect 65150 29696 65156 29708
rect 65015 29668 65156 29696
rect 65015 29665 65027 29668
rect 64969 29659 65027 29665
rect 65150 29656 65156 29668
rect 65208 29656 65214 29708
rect 65061 29631 65119 29637
rect 65061 29597 65073 29631
rect 65107 29628 65119 29631
rect 65889 29631 65947 29637
rect 65889 29628 65901 29631
rect 65107 29600 65901 29628
rect 65107 29597 65119 29600
rect 65061 29591 65119 29597
rect 65889 29597 65901 29600
rect 65935 29628 65947 29631
rect 66530 29628 66536 29640
rect 65935 29600 66536 29628
rect 65935 29597 65947 29600
rect 65889 29591 65947 29597
rect 66530 29588 66536 29600
rect 66588 29588 66594 29640
rect 64509 29495 64567 29501
rect 64509 29461 64521 29495
rect 64555 29492 64567 29495
rect 64690 29492 64696 29504
rect 64555 29464 64696 29492
rect 64555 29461 64567 29464
rect 64509 29455 64567 29461
rect 64690 29452 64696 29464
rect 64748 29452 64754 29504
rect 63572 29402 66424 29424
rect 63572 29350 64338 29402
rect 64390 29350 64402 29402
rect 64454 29350 64466 29402
rect 64518 29350 64530 29402
rect 64582 29350 64594 29402
rect 64646 29350 66424 29402
rect 63572 29328 66424 29350
rect 65610 29248 65616 29300
rect 65668 29288 65674 29300
rect 65797 29291 65855 29297
rect 65797 29288 65809 29291
rect 65668 29260 65809 29288
rect 65668 29248 65674 29260
rect 65797 29257 65809 29260
rect 65843 29257 65855 29291
rect 65797 29251 65855 29257
rect 64046 29112 64052 29164
rect 64104 29112 64110 29164
rect 64325 29155 64383 29161
rect 64325 29121 64337 29155
rect 64371 29152 64383 29155
rect 64690 29152 64696 29164
rect 64371 29124 64696 29152
rect 64371 29121 64383 29124
rect 64325 29115 64383 29121
rect 64690 29112 64696 29124
rect 64748 29112 64754 29164
rect 65794 29016 65800 29028
rect 65550 28988 65800 29016
rect 65794 28976 65800 28988
rect 65852 29016 65858 29028
rect 66438 29016 66444 29028
rect 65852 28988 66444 29016
rect 65852 28976 65858 28988
rect 66438 28976 66444 28988
rect 66496 28976 66502 29028
rect 63572 28858 66424 28880
rect 63572 28806 65258 28858
rect 65310 28806 65322 28858
rect 65374 28806 65386 28858
rect 65438 28806 65450 28858
rect 65502 28806 65514 28858
rect 65566 28806 66424 28858
rect 63572 28784 66424 28806
rect 63310 28704 63316 28756
rect 63368 28744 63374 28756
rect 64785 28747 64843 28753
rect 64785 28744 64797 28747
rect 63368 28716 64797 28744
rect 63368 28704 63374 28716
rect 64785 28713 64797 28716
rect 64831 28713 64843 28747
rect 64785 28707 64843 28713
rect 65150 28704 65156 28756
rect 65208 28704 65214 28756
rect 65978 28744 65984 28756
rect 65536 28716 65984 28744
rect 64693 28679 64751 28685
rect 64693 28645 64705 28679
rect 64739 28676 64751 28679
rect 64739 28648 64874 28676
rect 64739 28645 64751 28648
rect 64693 28639 64751 28645
rect 64846 28608 64874 28648
rect 65058 28636 65064 28688
rect 65116 28676 65122 28688
rect 65429 28679 65487 28685
rect 65429 28676 65441 28679
rect 65116 28648 65441 28676
rect 65116 28636 65122 28648
rect 65429 28645 65441 28648
rect 65475 28645 65487 28679
rect 65429 28639 65487 28645
rect 65536 28608 65564 28716
rect 65978 28704 65984 28716
rect 66036 28704 66042 28756
rect 64846 28580 65564 28608
rect 65610 28568 65616 28620
rect 65668 28608 65674 28620
rect 65981 28611 66039 28617
rect 65981 28608 65993 28611
rect 65668 28580 65993 28608
rect 65668 28568 65674 28580
rect 65981 28577 65993 28580
rect 66027 28577 66039 28611
rect 65981 28571 66039 28577
rect 64601 28543 64659 28549
rect 64601 28509 64613 28543
rect 64647 28509 64659 28543
rect 64601 28503 64659 28509
rect 64616 28472 64644 28503
rect 64874 28472 64880 28484
rect 64616 28444 64880 28472
rect 64874 28432 64880 28444
rect 64932 28472 64938 28484
rect 65150 28472 65156 28484
rect 64932 28444 65156 28472
rect 64932 28432 64938 28444
rect 65150 28432 65156 28444
rect 65208 28432 65214 28484
rect 63572 28314 66424 28336
rect 63572 28262 64338 28314
rect 64390 28262 64402 28314
rect 64454 28262 64466 28314
rect 64518 28262 64530 28314
rect 64582 28262 64594 28314
rect 64646 28262 66424 28314
rect 63572 28240 66424 28262
rect 63310 28160 63316 28212
rect 63368 28200 63374 28212
rect 64417 28203 64475 28209
rect 64417 28200 64429 28203
rect 63368 28172 64429 28200
rect 63368 28160 63374 28172
rect 64417 28169 64429 28172
rect 64463 28169 64475 28203
rect 64417 28163 64475 28169
rect 63572 27770 66424 27792
rect 63572 27718 65258 27770
rect 65310 27718 65322 27770
rect 65374 27718 65386 27770
rect 65438 27718 65450 27770
rect 65502 27718 65514 27770
rect 65566 27718 66424 27770
rect 63572 27696 66424 27718
rect 65061 27659 65119 27665
rect 65061 27625 65073 27659
rect 65107 27656 65119 27659
rect 65610 27656 65616 27668
rect 65107 27628 65616 27656
rect 65107 27625 65119 27628
rect 65061 27619 65119 27625
rect 65610 27616 65616 27628
rect 65668 27616 65674 27668
rect 64874 27480 64880 27532
rect 64932 27520 64938 27532
rect 64969 27523 65027 27529
rect 64969 27520 64981 27523
rect 64932 27492 64981 27520
rect 64932 27480 64938 27492
rect 64969 27489 64981 27492
rect 65015 27489 65027 27523
rect 64969 27483 65027 27489
rect 65150 27412 65156 27464
rect 65208 27452 65214 27464
rect 65245 27455 65303 27461
rect 65245 27452 65257 27455
rect 65208 27424 65257 27452
rect 65208 27412 65214 27424
rect 65245 27421 65257 27424
rect 65291 27452 65303 27455
rect 65702 27452 65708 27464
rect 65291 27424 65708 27452
rect 65291 27421 65303 27424
rect 65245 27415 65303 27421
rect 65702 27412 65708 27424
rect 65760 27412 65766 27464
rect 64601 27319 64659 27325
rect 64601 27285 64613 27319
rect 64647 27316 64659 27319
rect 65058 27316 65064 27328
rect 64647 27288 65064 27316
rect 64647 27285 64659 27288
rect 64601 27279 64659 27285
rect 65058 27276 65064 27288
rect 65116 27276 65122 27328
rect 63572 27226 66424 27248
rect 63572 27174 64338 27226
rect 64390 27174 64402 27226
rect 64454 27174 64466 27226
rect 64518 27174 64530 27226
rect 64582 27174 64594 27226
rect 64646 27174 66424 27226
rect 63572 27152 66424 27174
rect 64049 26979 64107 26985
rect 64049 26945 64061 26979
rect 64095 26976 64107 26979
rect 64690 26976 64696 26988
rect 64095 26948 64696 26976
rect 64095 26945 64107 26948
rect 64049 26939 64107 26945
rect 64690 26936 64696 26948
rect 64748 26936 64754 26988
rect 65794 26908 65800 26920
rect 65458 26880 65800 26908
rect 65794 26868 65800 26880
rect 65852 26908 65858 26920
rect 65978 26908 65984 26920
rect 65852 26880 65984 26908
rect 65852 26868 65858 26880
rect 65978 26868 65984 26880
rect 66036 26868 66042 26920
rect 64325 26843 64383 26849
rect 64325 26809 64337 26843
rect 64371 26840 64383 26843
rect 64598 26840 64604 26852
rect 64371 26812 64604 26840
rect 64371 26809 64383 26812
rect 64325 26803 64383 26809
rect 64598 26800 64604 26812
rect 64656 26800 64662 26852
rect 65794 26732 65800 26784
rect 65852 26732 65858 26784
rect 63572 26682 66424 26704
rect 63572 26630 65258 26682
rect 65310 26630 65322 26682
rect 65374 26630 65386 26682
rect 65438 26630 65450 26682
rect 65502 26630 65514 26682
rect 65566 26630 66424 26682
rect 63572 26608 66424 26630
rect 64598 26528 64604 26580
rect 64656 26528 64662 26580
rect 65058 26528 65064 26580
rect 65116 26528 65122 26580
rect 65518 26528 65524 26580
rect 65576 26568 65582 26580
rect 65978 26568 65984 26580
rect 65576 26540 65984 26568
rect 65576 26528 65582 26540
rect 65978 26528 65984 26540
rect 66036 26528 66042 26580
rect 64969 26435 65027 26441
rect 64969 26401 64981 26435
rect 65015 26432 65027 26435
rect 65429 26435 65487 26441
rect 65429 26432 65441 26435
rect 65015 26404 65441 26432
rect 65015 26401 65027 26404
rect 64969 26395 65027 26401
rect 65429 26401 65441 26404
rect 65475 26401 65487 26435
rect 65429 26395 65487 26401
rect 65794 26392 65800 26444
rect 65852 26432 65858 26444
rect 65978 26432 65984 26444
rect 65852 26404 65984 26432
rect 65852 26392 65858 26404
rect 65978 26392 65984 26404
rect 66036 26392 66042 26444
rect 65150 26324 65156 26376
rect 65208 26364 65214 26376
rect 65245 26367 65303 26373
rect 65245 26364 65257 26367
rect 65208 26336 65257 26364
rect 65208 26324 65214 26336
rect 65245 26333 65257 26336
rect 65291 26364 65303 26367
rect 66530 26364 66536 26376
rect 65291 26336 66536 26364
rect 65291 26333 65303 26336
rect 65245 26327 65303 26333
rect 66530 26324 66536 26336
rect 66588 26324 66594 26376
rect 64874 26256 64880 26308
rect 64932 26296 64938 26308
rect 65794 26296 65800 26308
rect 64932 26268 65800 26296
rect 64932 26256 64938 26268
rect 65794 26256 65800 26268
rect 65852 26256 65858 26308
rect 63862 26188 63868 26240
rect 63920 26228 63926 26240
rect 64046 26228 64052 26240
rect 63920 26200 64052 26228
rect 63920 26188 63926 26200
rect 64046 26188 64052 26200
rect 64104 26188 64110 26240
rect 63572 26138 66424 26160
rect 63572 26086 64338 26138
rect 64390 26086 64402 26138
rect 64454 26086 64466 26138
rect 64518 26086 64530 26138
rect 64582 26086 64594 26138
rect 64646 26086 66424 26138
rect 63572 26064 66424 26086
rect 63572 25594 66424 25616
rect 63572 25542 65258 25594
rect 65310 25542 65322 25594
rect 65374 25542 65386 25594
rect 65438 25542 65450 25594
rect 65502 25542 65514 25594
rect 65566 25542 66424 25594
rect 63572 25520 66424 25542
rect 63954 25304 63960 25356
rect 64012 25304 64018 25356
rect 64969 25347 65027 25353
rect 64969 25313 64981 25347
rect 65015 25344 65027 25347
rect 65429 25347 65487 25353
rect 65429 25344 65441 25347
rect 65015 25316 65441 25344
rect 65015 25313 65027 25316
rect 64969 25307 65027 25313
rect 65429 25313 65441 25316
rect 65475 25313 65487 25347
rect 65429 25307 65487 25313
rect 65058 25236 65064 25288
rect 65116 25236 65122 25288
rect 65150 25236 65156 25288
rect 65208 25236 65214 25288
rect 65794 25236 65800 25288
rect 65852 25276 65858 25288
rect 65981 25279 66039 25285
rect 65981 25276 65993 25279
rect 65852 25248 65993 25276
rect 65852 25236 65858 25248
rect 65981 25245 65993 25248
rect 66027 25245 66039 25279
rect 65981 25239 66039 25245
rect 64230 25100 64236 25152
rect 64288 25140 64294 25152
rect 64601 25143 64659 25149
rect 64601 25140 64613 25143
rect 64288 25112 64613 25140
rect 64288 25100 64294 25112
rect 64601 25109 64613 25112
rect 64647 25109 64659 25143
rect 64601 25103 64659 25109
rect 63572 25050 66424 25072
rect 63572 24998 64338 25050
rect 64390 24998 64402 25050
rect 64454 24998 64466 25050
rect 64518 24998 64530 25050
rect 64582 24998 64594 25050
rect 64646 24998 66424 25050
rect 63572 24976 66424 24998
rect 63218 24828 63224 24880
rect 63276 24868 63282 24880
rect 63586 24868 63592 24880
rect 63276 24840 63592 24868
rect 63276 24828 63282 24840
rect 63586 24828 63592 24840
rect 63644 24828 63650 24880
rect 63865 24735 63923 24741
rect 63865 24701 63877 24735
rect 63911 24732 63923 24735
rect 64966 24732 64972 24744
rect 63911 24704 64972 24732
rect 63911 24701 63923 24704
rect 63865 24695 63923 24701
rect 64966 24692 64972 24704
rect 65024 24692 65030 24744
rect 63954 24556 63960 24608
rect 64012 24596 64018 24608
rect 65153 24599 65211 24605
rect 65153 24596 65165 24599
rect 64012 24568 65165 24596
rect 64012 24556 64018 24568
rect 65153 24565 65165 24568
rect 65199 24565 65211 24599
rect 65153 24559 65211 24565
rect 63572 24506 66424 24528
rect 63572 24454 65258 24506
rect 65310 24454 65322 24506
rect 65374 24454 65386 24506
rect 65438 24454 65450 24506
rect 65502 24454 65514 24506
rect 65566 24454 66424 24506
rect 63572 24432 66424 24454
rect 64690 24352 64696 24404
rect 64748 24392 64754 24404
rect 65153 24395 65211 24401
rect 65153 24392 65165 24395
rect 64748 24364 65165 24392
rect 64748 24352 64754 24364
rect 65153 24361 65165 24364
rect 65199 24361 65211 24395
rect 65153 24355 65211 24361
rect 63865 24327 63923 24333
rect 63865 24293 63877 24327
rect 63911 24324 63923 24327
rect 64046 24324 64052 24336
rect 63911 24296 64052 24324
rect 63911 24293 63923 24296
rect 63865 24287 63923 24293
rect 64046 24284 64052 24296
rect 64104 24284 64110 24336
rect 63572 23962 66424 23984
rect 63572 23910 64338 23962
rect 64390 23910 64402 23962
rect 64454 23910 64466 23962
rect 64518 23910 64530 23962
rect 64582 23910 64594 23962
rect 64646 23910 66424 23962
rect 63572 23888 66424 23910
rect 63954 23604 63960 23656
rect 64012 23644 64018 23656
rect 64049 23647 64107 23653
rect 64049 23644 64061 23647
rect 64012 23616 64061 23644
rect 64012 23604 64018 23616
rect 64049 23613 64061 23616
rect 64095 23613 64107 23647
rect 64049 23607 64107 23613
rect 64230 23536 64236 23588
rect 64288 23576 64294 23588
rect 64325 23579 64383 23585
rect 64325 23576 64337 23579
rect 64288 23548 64337 23576
rect 64288 23536 64294 23548
rect 64325 23545 64337 23548
rect 64371 23545 64383 23579
rect 65610 23576 65616 23588
rect 65550 23548 65616 23576
rect 64325 23539 64383 23545
rect 65610 23536 65616 23548
rect 65668 23536 65674 23588
rect 63034 23468 63040 23520
rect 63092 23508 63098 23520
rect 63862 23508 63868 23520
rect 63092 23480 63868 23508
rect 63092 23468 63098 23480
rect 63862 23468 63868 23480
rect 63920 23468 63926 23520
rect 65794 23468 65800 23520
rect 65852 23468 65858 23520
rect 63572 23418 66424 23440
rect 63572 23366 65258 23418
rect 65310 23366 65322 23418
rect 65374 23366 65386 23418
rect 65438 23366 65450 23418
rect 65502 23366 65514 23418
rect 65566 23366 66424 23418
rect 63572 23344 66424 23366
rect 65058 23264 65064 23316
rect 65116 23304 65122 23316
rect 65245 23307 65303 23313
rect 65245 23304 65257 23307
rect 65116 23276 65257 23304
rect 65116 23264 65122 23276
rect 65245 23273 65257 23276
rect 65291 23273 65303 23307
rect 65245 23267 65303 23273
rect 64785 23239 64843 23245
rect 64785 23205 64797 23239
rect 64831 23236 64843 23239
rect 65978 23236 65984 23248
rect 64831 23208 65984 23236
rect 64831 23205 64843 23208
rect 64785 23199 64843 23205
rect 65978 23196 65984 23208
rect 66036 23196 66042 23248
rect 64417 23171 64475 23177
rect 64417 23137 64429 23171
rect 64463 23168 64475 23171
rect 64874 23168 64880 23180
rect 64463 23140 64880 23168
rect 64463 23137 64475 23140
rect 64417 23131 64475 23137
rect 64874 23128 64880 23140
rect 64932 23168 64938 23180
rect 65886 23168 65892 23180
rect 64932 23140 65892 23168
rect 64932 23128 64938 23140
rect 65886 23128 65892 23140
rect 65944 23128 65950 23180
rect 64693 23103 64751 23109
rect 64693 23069 64705 23103
rect 64739 23100 64751 23103
rect 65702 23100 65708 23112
rect 64739 23072 65708 23100
rect 64739 23069 64751 23072
rect 64693 23063 64751 23069
rect 65702 23060 65708 23072
rect 65760 23060 65766 23112
rect 63572 22874 66424 22896
rect 63572 22822 64338 22874
rect 64390 22822 64402 22874
rect 64454 22822 64466 22874
rect 64518 22822 64530 22874
rect 64582 22822 64594 22874
rect 64646 22822 66424 22874
rect 63572 22800 66424 22822
rect 64601 22763 64659 22769
rect 64601 22729 64613 22763
rect 64647 22760 64659 22763
rect 64874 22760 64880 22772
rect 64647 22732 64880 22760
rect 64647 22729 64659 22732
rect 64601 22723 64659 22729
rect 64874 22720 64880 22732
rect 64932 22720 64938 22772
rect 64046 22516 64052 22568
rect 64104 22556 64110 22568
rect 64325 22559 64383 22565
rect 64325 22556 64337 22559
rect 64104 22528 64337 22556
rect 64104 22516 64110 22528
rect 64325 22525 64337 22528
rect 64371 22556 64383 22559
rect 64690 22556 64696 22568
rect 64371 22528 64696 22556
rect 64371 22525 64383 22528
rect 64325 22519 64383 22525
rect 64690 22516 64696 22528
rect 64748 22516 64754 22568
rect 64138 22448 64144 22500
rect 64196 22488 64202 22500
rect 64874 22488 64880 22500
rect 64196 22460 64880 22488
rect 64196 22448 64202 22460
rect 64874 22448 64880 22460
rect 64932 22488 64938 22500
rect 65337 22491 65395 22497
rect 65337 22488 65349 22491
rect 64932 22460 65349 22488
rect 64932 22448 64938 22460
rect 65337 22457 65349 22460
rect 65383 22457 65395 22491
rect 65337 22451 65395 22457
rect 65705 22491 65763 22497
rect 65705 22457 65717 22491
rect 65751 22488 65763 22491
rect 65886 22488 65892 22500
rect 65751 22460 65892 22488
rect 65751 22457 65763 22460
rect 65705 22451 65763 22457
rect 65886 22448 65892 22460
rect 65944 22448 65950 22500
rect 63572 22330 66424 22352
rect 63572 22278 65258 22330
rect 65310 22278 65322 22330
rect 65374 22278 65386 22330
rect 65438 22278 65450 22330
rect 65502 22278 65514 22330
rect 65566 22278 66424 22330
rect 63572 22256 66424 22278
rect 65797 22219 65855 22225
rect 65797 22185 65809 22219
rect 65843 22216 65855 22219
rect 66254 22216 66260 22228
rect 65843 22188 66260 22216
rect 65843 22185 65855 22188
rect 65797 22179 65855 22185
rect 66254 22176 66260 22188
rect 66312 22176 66318 22228
rect 65886 22148 65892 22160
rect 65550 22120 65892 22148
rect 65886 22108 65892 22120
rect 65944 22108 65950 22160
rect 63954 22040 63960 22092
rect 64012 22080 64018 22092
rect 64049 22083 64107 22089
rect 64049 22080 64061 22083
rect 64012 22052 64061 22080
rect 64012 22040 64018 22052
rect 64049 22049 64061 22052
rect 64095 22049 64107 22083
rect 64049 22043 64107 22049
rect 64325 22015 64383 22021
rect 64325 21981 64337 22015
rect 64371 22012 64383 22015
rect 64690 22012 64696 22024
rect 64371 21984 64696 22012
rect 64371 21981 64383 21984
rect 64325 21975 64383 21981
rect 64690 21972 64696 21984
rect 64748 21972 64754 22024
rect 63572 21786 66424 21808
rect 63572 21734 64338 21786
rect 64390 21734 64402 21786
rect 64454 21734 64466 21786
rect 64518 21734 64530 21786
rect 64582 21734 64594 21786
rect 64646 21734 66424 21786
rect 63572 21712 66424 21734
rect 65702 21428 65708 21480
rect 65760 21468 65766 21480
rect 65981 21471 66039 21477
rect 65981 21468 65993 21471
rect 65760 21440 65993 21468
rect 65760 21428 65766 21440
rect 65981 21437 65993 21440
rect 66027 21468 66039 21471
rect 66254 21468 66260 21480
rect 66027 21440 66260 21468
rect 66027 21437 66039 21440
rect 65981 21431 66039 21437
rect 66254 21428 66260 21440
rect 66312 21428 66318 21480
rect 63310 21360 63316 21412
rect 63368 21400 63374 21412
rect 63862 21400 63868 21412
rect 63368 21372 63868 21400
rect 63368 21360 63374 21372
rect 63862 21360 63868 21372
rect 63920 21400 63926 21412
rect 64969 21403 65027 21409
rect 64969 21400 64981 21403
rect 63920 21372 64981 21400
rect 63920 21360 63926 21372
rect 64969 21369 64981 21372
rect 65015 21369 65027 21403
rect 64969 21363 65027 21369
rect 65337 21403 65395 21409
rect 65337 21369 65349 21403
rect 65383 21400 65395 21403
rect 65610 21400 65616 21412
rect 65383 21372 65616 21400
rect 65383 21369 65395 21372
rect 65337 21363 65395 21369
rect 65610 21360 65616 21372
rect 65668 21360 65674 21412
rect 65150 21292 65156 21344
rect 65208 21332 65214 21344
rect 65429 21335 65487 21341
rect 65429 21332 65441 21335
rect 65208 21304 65441 21332
rect 65208 21292 65214 21304
rect 65429 21301 65441 21304
rect 65475 21301 65487 21335
rect 65429 21295 65487 21301
rect 63572 21242 66424 21264
rect 63572 21190 65258 21242
rect 65310 21190 65322 21242
rect 65374 21190 65386 21242
rect 65438 21190 65450 21242
rect 65502 21190 65514 21242
rect 65566 21190 66424 21242
rect 63572 21168 66424 21190
rect 64601 21131 64659 21137
rect 64601 21097 64613 21131
rect 64647 21128 64659 21131
rect 64690 21128 64696 21140
rect 64647 21100 64696 21128
rect 64647 21097 64659 21100
rect 64601 21091 64659 21097
rect 64690 21088 64696 21100
rect 64748 21088 64754 21140
rect 64969 21131 65027 21137
rect 64969 21097 64981 21131
rect 65015 21128 65027 21131
rect 65150 21128 65156 21140
rect 65015 21100 65156 21128
rect 65015 21097 65027 21100
rect 64969 21091 65027 21097
rect 65150 21088 65156 21100
rect 65208 21088 65214 21140
rect 65058 20884 65064 20936
rect 65116 20884 65122 20936
rect 65245 20927 65303 20933
rect 65245 20893 65257 20927
rect 65291 20924 65303 20927
rect 65610 20924 65616 20936
rect 65291 20896 65616 20924
rect 65291 20893 65303 20896
rect 65245 20887 65303 20893
rect 65610 20884 65616 20896
rect 65668 20884 65674 20936
rect 63572 20698 66424 20720
rect 63572 20646 64338 20698
rect 64390 20646 64402 20698
rect 64454 20646 64466 20698
rect 64518 20646 64530 20698
rect 64582 20646 64594 20698
rect 64646 20646 66424 20698
rect 63572 20624 66424 20646
rect 64966 20408 64972 20460
rect 65024 20448 65030 20460
rect 65153 20451 65211 20457
rect 65153 20448 65165 20451
rect 65024 20420 65165 20448
rect 65024 20408 65030 20420
rect 65153 20417 65165 20420
rect 65199 20417 65211 20451
rect 65153 20411 65211 20417
rect 65061 20383 65119 20389
rect 65061 20349 65073 20383
rect 65107 20380 65119 20383
rect 65794 20380 65800 20392
rect 65107 20352 65800 20380
rect 65107 20349 65119 20352
rect 65061 20343 65119 20349
rect 65794 20340 65800 20352
rect 65852 20340 65858 20392
rect 64138 20272 64144 20324
rect 64196 20312 64202 20324
rect 66162 20312 66168 20324
rect 64196 20284 66168 20312
rect 64196 20272 64202 20284
rect 66162 20272 66168 20284
rect 66220 20272 66226 20324
rect 64601 20247 64659 20253
rect 64601 20213 64613 20247
rect 64647 20244 64659 20247
rect 64874 20244 64880 20256
rect 64647 20216 64880 20244
rect 64647 20213 64659 20216
rect 64601 20207 64659 20213
rect 64874 20204 64880 20216
rect 64932 20204 64938 20256
rect 64969 20247 65027 20253
rect 64969 20213 64981 20247
rect 65015 20244 65027 20247
rect 65794 20244 65800 20256
rect 65015 20216 65800 20244
rect 65015 20213 65027 20216
rect 64969 20207 65027 20213
rect 65794 20204 65800 20216
rect 65852 20204 65858 20256
rect 63572 20154 66424 20176
rect 63572 20102 65258 20154
rect 65310 20102 65322 20154
rect 65374 20102 65386 20154
rect 65438 20102 65450 20154
rect 65502 20102 65514 20154
rect 65566 20102 66424 20154
rect 63572 20080 66424 20102
rect 65886 19972 65892 19984
rect 65550 19944 65892 19972
rect 65886 19932 65892 19944
rect 65944 19972 65950 19984
rect 66162 19972 66168 19984
rect 65944 19944 66168 19972
rect 65944 19932 65950 19944
rect 66162 19932 66168 19944
rect 66220 19932 66226 19984
rect 64046 19796 64052 19848
rect 64104 19796 64110 19848
rect 64325 19839 64383 19845
rect 64325 19805 64337 19839
rect 64371 19836 64383 19839
rect 64690 19836 64696 19848
rect 64371 19808 64696 19836
rect 64371 19805 64383 19808
rect 64325 19799 64383 19805
rect 64690 19796 64696 19808
rect 64748 19796 64754 19848
rect 65797 19703 65855 19709
rect 65797 19669 65809 19703
rect 65843 19700 65855 19703
rect 65886 19700 65892 19712
rect 65843 19672 65892 19700
rect 65843 19669 65855 19672
rect 65797 19663 65855 19669
rect 65886 19660 65892 19672
rect 65944 19660 65950 19712
rect 63572 19610 66424 19632
rect 63572 19558 64338 19610
rect 64390 19558 64402 19610
rect 64454 19558 64466 19610
rect 64518 19558 64530 19610
rect 64582 19558 64594 19610
rect 64646 19558 66424 19610
rect 63572 19536 66424 19558
rect 64601 19499 64659 19505
rect 64601 19465 64613 19499
rect 64647 19496 64659 19499
rect 64690 19496 64696 19508
rect 64647 19468 64696 19496
rect 64647 19465 64659 19468
rect 64601 19459 64659 19465
rect 64690 19456 64696 19468
rect 64748 19456 64754 19508
rect 65245 19363 65303 19369
rect 65245 19329 65257 19363
rect 65291 19360 65303 19363
rect 65610 19360 65616 19372
rect 65291 19332 65616 19360
rect 65291 19329 65303 19332
rect 65245 19323 65303 19329
rect 65610 19320 65616 19332
rect 65668 19320 65674 19372
rect 64874 19252 64880 19304
rect 64932 19292 64938 19304
rect 65061 19295 65119 19301
rect 65061 19292 65073 19295
rect 64932 19264 65073 19292
rect 64932 19252 64938 19264
rect 65061 19261 65073 19264
rect 65107 19261 65119 19295
rect 65061 19255 65119 19261
rect 65886 19252 65892 19304
rect 65944 19292 65950 19304
rect 65981 19295 66039 19301
rect 65981 19292 65993 19295
rect 65944 19264 65993 19292
rect 65944 19252 65950 19264
rect 65981 19261 65993 19264
rect 66027 19261 66039 19295
rect 65981 19255 66039 19261
rect 64969 19227 65027 19233
rect 64969 19193 64981 19227
rect 65015 19224 65027 19227
rect 65429 19227 65487 19233
rect 65429 19224 65441 19227
rect 65015 19196 65441 19224
rect 65015 19193 65027 19196
rect 64969 19187 65027 19193
rect 65429 19193 65441 19196
rect 65475 19193 65487 19227
rect 65429 19187 65487 19193
rect 63572 19066 66424 19088
rect 63572 19014 65258 19066
rect 65310 19014 65322 19066
rect 65374 19014 65386 19066
rect 65438 19014 65450 19066
rect 65502 19014 65514 19066
rect 65566 19014 66424 19066
rect 63572 18992 66424 19014
rect 64969 18819 65027 18825
rect 64969 18785 64981 18819
rect 65015 18816 65027 18819
rect 65429 18819 65487 18825
rect 65429 18816 65441 18819
rect 65015 18788 65441 18816
rect 65015 18785 65027 18788
rect 64969 18779 65027 18785
rect 65429 18785 65441 18788
rect 65475 18785 65487 18819
rect 65429 18779 65487 18785
rect 65058 18708 65064 18760
rect 65116 18708 65122 18760
rect 65245 18751 65303 18757
rect 65245 18717 65257 18751
rect 65291 18748 65303 18751
rect 65610 18748 65616 18760
rect 65291 18720 65616 18748
rect 65291 18717 65303 18720
rect 65245 18711 65303 18717
rect 65610 18708 65616 18720
rect 65668 18708 65674 18760
rect 65978 18708 65984 18760
rect 66036 18708 66042 18760
rect 64601 18615 64659 18621
rect 64601 18581 64613 18615
rect 64647 18612 64659 18615
rect 64690 18612 64696 18624
rect 64647 18584 64696 18612
rect 64647 18581 64659 18584
rect 64601 18575 64659 18581
rect 64690 18572 64696 18584
rect 64748 18572 64754 18624
rect 63572 18522 66424 18544
rect 63572 18470 64338 18522
rect 64390 18470 64402 18522
rect 64454 18470 64466 18522
rect 64518 18470 64530 18522
rect 64582 18470 64594 18522
rect 64646 18470 66424 18522
rect 63572 18448 66424 18470
rect 63034 18368 63040 18420
rect 63092 18408 63098 18420
rect 66070 18408 66076 18420
rect 63092 18380 66076 18408
rect 63092 18368 63098 18380
rect 66070 18368 66076 18380
rect 66128 18368 66134 18420
rect 64325 18275 64383 18281
rect 64325 18241 64337 18275
rect 64371 18272 64383 18275
rect 64690 18272 64696 18284
rect 64371 18244 64696 18272
rect 64371 18241 64383 18244
rect 64325 18235 64383 18241
rect 64690 18232 64696 18244
rect 64748 18232 64754 18284
rect 64046 18164 64052 18216
rect 64104 18164 64110 18216
rect 66162 18136 66168 18148
rect 65550 18108 66168 18136
rect 66162 18096 66168 18108
rect 66220 18096 66226 18148
rect 64966 18028 64972 18080
rect 65024 18068 65030 18080
rect 65797 18071 65855 18077
rect 65797 18068 65809 18071
rect 65024 18040 65809 18068
rect 65024 18028 65030 18040
rect 65797 18037 65809 18040
rect 65843 18068 65855 18071
rect 65978 18068 65984 18080
rect 65843 18040 65984 18068
rect 65843 18037 65855 18040
rect 65797 18031 65855 18037
rect 65978 18028 65984 18040
rect 66036 18028 66042 18080
rect 63572 17978 66424 18000
rect 63572 17926 65258 17978
rect 65310 17926 65322 17978
rect 65374 17926 65386 17978
rect 65438 17926 65450 17978
rect 65502 17926 65514 17978
rect 65566 17926 66424 17978
rect 63572 17904 66424 17926
rect 64785 17867 64843 17873
rect 64785 17833 64797 17867
rect 64831 17864 64843 17867
rect 64966 17864 64972 17876
rect 64831 17836 64972 17864
rect 64831 17833 64843 17836
rect 64785 17827 64843 17833
rect 64966 17824 64972 17836
rect 65024 17824 65030 17876
rect 65058 17824 65064 17876
rect 65116 17864 65122 17876
rect 65337 17867 65395 17873
rect 65337 17864 65349 17867
rect 65116 17836 65349 17864
rect 65116 17824 65122 17836
rect 65337 17833 65349 17836
rect 65383 17833 65395 17867
rect 65337 17827 65395 17833
rect 65702 17824 65708 17876
rect 65760 17824 65766 17876
rect 64690 17756 64696 17808
rect 64748 17796 64754 17808
rect 64877 17799 64935 17805
rect 64877 17796 64889 17799
rect 64748 17768 64889 17796
rect 64748 17756 64754 17768
rect 64877 17765 64889 17768
rect 64923 17765 64935 17799
rect 64877 17759 64935 17765
rect 65797 17731 65855 17737
rect 65797 17697 65809 17731
rect 65843 17728 65855 17731
rect 65978 17728 65984 17740
rect 65843 17700 65984 17728
rect 65843 17697 65855 17700
rect 65797 17691 65855 17697
rect 65978 17688 65984 17700
rect 66036 17688 66042 17740
rect 64693 17663 64751 17669
rect 64693 17629 64705 17663
rect 64739 17660 64751 17663
rect 64874 17660 64880 17672
rect 64739 17632 64880 17660
rect 64739 17629 64751 17632
rect 64693 17623 64751 17629
rect 64874 17620 64880 17632
rect 64932 17660 64938 17672
rect 65889 17663 65947 17669
rect 65889 17660 65901 17663
rect 64932 17632 65901 17660
rect 64932 17620 64938 17632
rect 65889 17629 65901 17632
rect 65935 17629 65947 17663
rect 65889 17623 65947 17629
rect 65150 17552 65156 17604
rect 65208 17592 65214 17604
rect 65245 17595 65303 17601
rect 65245 17592 65257 17595
rect 65208 17564 65257 17592
rect 65208 17552 65214 17564
rect 65245 17561 65257 17564
rect 65291 17561 65303 17595
rect 65245 17555 65303 17561
rect 63572 17434 66424 17456
rect 63572 17382 64338 17434
rect 64390 17382 64402 17434
rect 64454 17382 64466 17434
rect 64518 17382 64530 17434
rect 64582 17382 64594 17434
rect 64646 17382 66424 17434
rect 63572 17360 66424 17382
rect 64601 17323 64659 17329
rect 64601 17289 64613 17323
rect 64647 17320 64659 17323
rect 64690 17320 64696 17332
rect 64647 17292 64696 17320
rect 64647 17289 64659 17292
rect 64601 17283 64659 17289
rect 64690 17280 64696 17292
rect 64748 17280 64754 17332
rect 63572 16890 66424 16912
rect 63572 16838 65258 16890
rect 65310 16838 65322 16890
rect 65374 16838 65386 16890
rect 65438 16838 65450 16890
rect 65502 16838 65514 16890
rect 65566 16838 66424 16890
rect 63572 16816 66424 16838
rect 62942 16668 62948 16720
rect 63000 16708 63006 16720
rect 66070 16708 66076 16720
rect 63000 16680 66076 16708
rect 63000 16668 63006 16680
rect 66070 16668 66076 16680
rect 66128 16668 66134 16720
rect 63310 16600 63316 16652
rect 63368 16600 63374 16652
rect 64969 16643 65027 16649
rect 64969 16609 64981 16643
rect 65015 16640 65027 16643
rect 65429 16643 65487 16649
rect 65429 16640 65441 16643
rect 65015 16612 65441 16640
rect 65015 16609 65027 16612
rect 64969 16603 65027 16609
rect 65429 16609 65441 16612
rect 65475 16609 65487 16643
rect 65429 16603 65487 16609
rect 65794 16600 65800 16652
rect 65852 16640 65858 16652
rect 65981 16643 66039 16649
rect 65981 16640 65993 16643
rect 65852 16612 65993 16640
rect 65852 16600 65858 16612
rect 65981 16609 65993 16612
rect 66027 16609 66039 16643
rect 65981 16603 66039 16609
rect 63328 16572 63356 16600
rect 63328 16544 63540 16572
rect 63512 16504 63540 16544
rect 65058 16532 65064 16584
rect 65116 16532 65122 16584
rect 65153 16575 65211 16581
rect 65153 16541 65165 16575
rect 65199 16541 65211 16575
rect 65153 16535 65211 16541
rect 65168 16504 65196 16535
rect 63512 16476 65196 16504
rect 63512 16448 63540 16476
rect 63494 16396 63500 16448
rect 63552 16396 63558 16448
rect 64601 16439 64659 16445
rect 64601 16405 64613 16439
rect 64647 16436 64659 16439
rect 64690 16436 64696 16448
rect 64647 16408 64696 16436
rect 64647 16405 64659 16408
rect 64601 16399 64659 16405
rect 64690 16396 64696 16408
rect 64748 16396 64754 16448
rect 63572 16346 66424 16368
rect 63572 16294 64338 16346
rect 64390 16294 64402 16346
rect 64454 16294 64466 16346
rect 64518 16294 64530 16346
rect 64582 16294 64594 16346
rect 64646 16294 66424 16346
rect 63572 16272 66424 16294
rect 65794 16192 65800 16244
rect 65852 16192 65858 16244
rect 63954 16056 63960 16108
rect 64012 16096 64018 16108
rect 64049 16099 64107 16105
rect 64049 16096 64061 16099
rect 64012 16068 64061 16096
rect 64012 16056 64018 16068
rect 64049 16065 64061 16068
rect 64095 16065 64107 16099
rect 64049 16059 64107 16065
rect 64325 16099 64383 16105
rect 64325 16065 64337 16099
rect 64371 16096 64383 16099
rect 64690 16096 64696 16108
rect 64371 16068 64696 16096
rect 64371 16065 64383 16068
rect 64325 16059 64383 16065
rect 64690 16056 64696 16068
rect 64748 16056 64754 16108
rect 66162 15960 66168 15972
rect 65550 15932 66168 15960
rect 66162 15920 66168 15932
rect 66220 15920 66226 15972
rect 63572 15802 66424 15824
rect 63572 15750 65258 15802
rect 65310 15750 65322 15802
rect 65374 15750 65386 15802
rect 65438 15750 65450 15802
rect 65502 15750 65514 15802
rect 65566 15750 66424 15802
rect 63572 15728 66424 15750
rect 64782 15648 64788 15700
rect 64840 15688 64846 15700
rect 64969 15691 65027 15697
rect 64969 15688 64981 15691
rect 64840 15660 64981 15688
rect 64840 15648 64846 15660
rect 64969 15657 64981 15660
rect 65015 15657 65027 15691
rect 64969 15651 65027 15657
rect 65058 15648 65064 15700
rect 65116 15688 65122 15700
rect 65337 15691 65395 15697
rect 65337 15688 65349 15691
rect 65116 15660 65349 15688
rect 65116 15648 65122 15660
rect 65337 15657 65349 15660
rect 65383 15657 65395 15691
rect 65337 15651 65395 15657
rect 64877 15623 64935 15629
rect 64877 15589 64889 15623
rect 64923 15620 64935 15623
rect 65886 15620 65892 15632
rect 64923 15592 65892 15620
rect 64923 15589 64935 15592
rect 64877 15583 64935 15589
rect 65886 15580 65892 15592
rect 65944 15580 65950 15632
rect 64785 15487 64843 15493
rect 64785 15453 64797 15487
rect 64831 15484 64843 15487
rect 64874 15484 64880 15496
rect 64831 15456 64880 15484
rect 64831 15453 64843 15456
rect 64785 15447 64843 15453
rect 64874 15444 64880 15456
rect 64932 15484 64938 15496
rect 65150 15484 65156 15496
rect 64932 15456 65156 15484
rect 64932 15444 64938 15456
rect 65150 15444 65156 15456
rect 65208 15444 65214 15496
rect 63572 15258 66424 15280
rect 63572 15206 64338 15258
rect 64390 15206 64402 15258
rect 64454 15206 64466 15258
rect 64518 15206 64530 15258
rect 64582 15206 64594 15258
rect 64646 15206 66424 15258
rect 63572 15184 66424 15206
rect 64693 15147 64751 15153
rect 64693 15113 64705 15147
rect 64739 15144 64751 15147
rect 64782 15144 64788 15156
rect 64739 15116 64788 15144
rect 64739 15113 64751 15116
rect 64693 15107 64751 15113
rect 64782 15104 64788 15116
rect 64840 15104 64846 15156
rect 63572 14714 66424 14736
rect 63572 14662 65258 14714
rect 65310 14662 65322 14714
rect 65374 14662 65386 14714
rect 65438 14662 65450 14714
rect 65502 14662 65514 14714
rect 65566 14662 66424 14714
rect 63572 14640 66424 14662
rect 63572 14170 66424 14192
rect 63572 14118 64338 14170
rect 64390 14118 64402 14170
rect 64454 14118 64466 14170
rect 64518 14118 64530 14170
rect 64582 14118 64594 14170
rect 64646 14118 66424 14170
rect 63572 14096 66424 14118
rect 63572 13626 66424 13648
rect 63572 13574 65258 13626
rect 65310 13574 65322 13626
rect 65374 13574 65386 13626
rect 65438 13574 65450 13626
rect 65502 13574 65514 13626
rect 65566 13574 66424 13626
rect 63572 13552 66424 13574
rect 63572 13082 66424 13104
rect 63572 13030 64338 13082
rect 64390 13030 64402 13082
rect 64454 13030 64466 13082
rect 64518 13030 64530 13082
rect 64582 13030 64594 13082
rect 64646 13030 66424 13082
rect 63572 13008 66424 13030
rect 63954 12792 63960 12844
rect 64012 12832 64018 12844
rect 64049 12835 64107 12841
rect 64049 12832 64061 12835
rect 64012 12804 64061 12832
rect 64012 12792 64018 12804
rect 64049 12801 64061 12804
rect 64095 12801 64107 12835
rect 64049 12795 64107 12801
rect 64325 12835 64383 12841
rect 64325 12801 64337 12835
rect 64371 12832 64383 12835
rect 65058 12832 65064 12844
rect 64371 12804 65064 12832
rect 64371 12801 64383 12804
rect 64325 12795 64383 12801
rect 65058 12792 65064 12804
rect 65116 12792 65122 12844
rect 66070 12792 66076 12844
rect 66128 12792 66134 12844
rect 64782 12696 64788 12708
rect 64708 12668 64788 12696
rect 64708 12628 64736 12668
rect 64782 12656 64788 12668
rect 64840 12656 64846 12708
rect 66438 12628 66444 12640
rect 64708 12600 66444 12628
rect 66438 12588 66444 12600
rect 66496 12588 66502 12640
rect 63572 12538 66424 12560
rect 63572 12486 65258 12538
rect 65310 12486 65322 12538
rect 65374 12486 65386 12538
rect 65438 12486 65450 12538
rect 65502 12486 65514 12538
rect 65566 12486 66424 12538
rect 63572 12464 66424 12486
rect 65797 12427 65855 12433
rect 65797 12393 65809 12427
rect 65843 12424 65855 12427
rect 65978 12424 65984 12436
rect 65843 12396 65984 12424
rect 65843 12393 65855 12396
rect 65797 12387 65855 12393
rect 65978 12384 65984 12396
rect 66036 12384 66042 12436
rect 66162 12356 66168 12368
rect 65550 12328 66168 12356
rect 66162 12316 66168 12328
rect 66220 12316 66226 12368
rect 63862 12180 63868 12232
rect 63920 12220 63926 12232
rect 64049 12223 64107 12229
rect 64049 12220 64061 12223
rect 63920 12192 64061 12220
rect 63920 12180 63926 12192
rect 64049 12189 64061 12192
rect 64095 12189 64107 12223
rect 64049 12183 64107 12189
rect 64325 12223 64383 12229
rect 64325 12189 64337 12223
rect 64371 12220 64383 12223
rect 64690 12220 64696 12232
rect 64371 12192 64696 12220
rect 64371 12189 64383 12192
rect 64325 12183 64383 12189
rect 64690 12180 64696 12192
rect 64748 12180 64754 12232
rect 63572 11994 66424 12016
rect 63572 11942 64338 11994
rect 64390 11942 64402 11994
rect 64454 11942 64466 11994
rect 64518 11942 64530 11994
rect 64582 11942 64594 11994
rect 64646 11942 66424 11994
rect 63572 11920 66424 11942
rect 64509 11883 64567 11889
rect 64509 11849 64521 11883
rect 64555 11880 64567 11883
rect 64690 11880 64696 11892
rect 64555 11852 64696 11880
rect 64555 11849 64567 11852
rect 64509 11843 64567 11849
rect 64690 11840 64696 11852
rect 64748 11840 64754 11892
rect 65058 11840 65064 11892
rect 65116 11880 65122 11892
rect 65337 11883 65395 11889
rect 65337 11880 65349 11883
rect 65116 11852 65349 11880
rect 65116 11840 65122 11852
rect 65337 11849 65349 11852
rect 65383 11849 65395 11883
rect 65337 11843 65395 11849
rect 65153 11747 65211 11753
rect 65153 11713 65165 11747
rect 65199 11744 65211 11747
rect 65610 11744 65616 11756
rect 65199 11716 65616 11744
rect 65199 11713 65211 11716
rect 65153 11707 65211 11713
rect 65610 11704 65616 11716
rect 65668 11744 65674 11756
rect 65889 11747 65947 11753
rect 65889 11744 65901 11747
rect 65668 11716 65901 11744
rect 65668 11704 65674 11716
rect 65889 11713 65901 11716
rect 65935 11713 65947 11747
rect 65889 11707 65947 11713
rect 62942 11636 62948 11688
rect 63000 11676 63006 11688
rect 64138 11676 64144 11688
rect 63000 11648 64144 11676
rect 63000 11636 63006 11648
rect 64138 11636 64144 11648
rect 64196 11636 64202 11688
rect 64969 11679 65027 11685
rect 64969 11645 64981 11679
rect 65015 11676 65027 11679
rect 66254 11676 66260 11688
rect 65015 11648 66260 11676
rect 65015 11645 65027 11648
rect 64969 11639 65027 11645
rect 66254 11636 66260 11648
rect 66312 11636 66318 11688
rect 65705 11611 65763 11617
rect 65705 11577 65717 11611
rect 65751 11608 65763 11611
rect 66070 11608 66076 11620
rect 65751 11580 66076 11608
rect 65751 11577 65763 11580
rect 65705 11571 65763 11577
rect 66070 11568 66076 11580
rect 66128 11568 66134 11620
rect 64874 11500 64880 11552
rect 64932 11500 64938 11552
rect 65797 11543 65855 11549
rect 65797 11509 65809 11543
rect 65843 11540 65855 11543
rect 65886 11540 65892 11552
rect 65843 11512 65892 11540
rect 65843 11509 65855 11512
rect 65797 11503 65855 11509
rect 65886 11500 65892 11512
rect 65944 11500 65950 11552
rect 63572 11450 66424 11472
rect 63572 11398 65258 11450
rect 65310 11398 65322 11450
rect 65374 11398 65386 11450
rect 65438 11398 65450 11450
rect 65502 11398 65514 11450
rect 65566 11398 66424 11450
rect 63572 11376 66424 11398
rect 64874 11296 64880 11348
rect 64932 11336 64938 11348
rect 65429 11339 65487 11345
rect 65429 11336 65441 11339
rect 64932 11308 65441 11336
rect 64932 11296 64938 11308
rect 65429 11305 65441 11308
rect 65475 11305 65487 11339
rect 65429 11299 65487 11305
rect 65978 11160 65984 11212
rect 66036 11160 66042 11212
rect 63572 10906 66424 10928
rect 63572 10854 64338 10906
rect 64390 10854 64402 10906
rect 64454 10854 64466 10906
rect 64518 10854 64530 10906
rect 64582 10854 64594 10906
rect 64646 10854 66424 10906
rect 63572 10832 66424 10854
rect 64601 10727 64659 10733
rect 64601 10693 64613 10727
rect 64647 10724 64659 10727
rect 65610 10724 65616 10736
rect 64647 10696 65616 10724
rect 64647 10693 64659 10696
rect 64601 10687 64659 10693
rect 65610 10684 65616 10696
rect 65668 10684 65674 10736
rect 65150 10616 65156 10668
rect 65208 10616 65214 10668
rect 65061 10591 65119 10597
rect 65061 10557 65073 10591
rect 65107 10588 65119 10591
rect 65794 10588 65800 10600
rect 65107 10560 65800 10588
rect 65107 10557 65119 10560
rect 65061 10551 65119 10557
rect 65794 10548 65800 10560
rect 65852 10548 65858 10600
rect 64966 10412 64972 10464
rect 65024 10412 65030 10464
rect 63572 10362 66424 10384
rect 63572 10310 65258 10362
rect 65310 10310 65322 10362
rect 65374 10310 65386 10362
rect 65438 10310 65450 10362
rect 65502 10310 65514 10362
rect 65566 10310 66424 10362
rect 63572 10288 66424 10310
rect 66162 10180 66168 10192
rect 65550 10152 66168 10180
rect 66162 10140 66168 10152
rect 66220 10140 66226 10192
rect 63862 10004 63868 10056
rect 63920 10044 63926 10056
rect 64049 10047 64107 10053
rect 64049 10044 64061 10047
rect 63920 10016 64061 10044
rect 63920 10004 63926 10016
rect 64049 10013 64061 10016
rect 64095 10013 64107 10047
rect 64049 10007 64107 10013
rect 64325 10047 64383 10053
rect 64325 10013 64337 10047
rect 64371 10044 64383 10047
rect 64690 10044 64696 10056
rect 64371 10016 64696 10044
rect 64371 10013 64383 10016
rect 64325 10007 64383 10013
rect 64690 10004 64696 10016
rect 64748 10004 64754 10056
rect 64966 9868 64972 9920
rect 65024 9908 65030 9920
rect 65797 9911 65855 9917
rect 65797 9908 65809 9911
rect 65024 9880 65809 9908
rect 65024 9868 65030 9880
rect 65797 9877 65809 9880
rect 65843 9877 65855 9911
rect 65797 9871 65855 9877
rect 63572 9818 66424 9840
rect 63572 9766 64338 9818
rect 64390 9766 64402 9818
rect 64454 9766 64466 9818
rect 64518 9766 64530 9818
rect 64582 9766 64594 9818
rect 64646 9766 66424 9818
rect 63572 9744 66424 9766
rect 63218 9596 63224 9648
rect 63276 9636 63282 9648
rect 63954 9636 63960 9648
rect 63276 9608 63960 9636
rect 63276 9596 63282 9608
rect 63954 9596 63960 9608
rect 64012 9596 64018 9648
rect 64800 9608 65056 9636
rect 64800 9500 64828 9608
rect 65028 9568 65056 9608
rect 65150 9568 65156 9580
rect 65208 9577 65214 9580
rect 65208 9571 65237 9577
rect 65028 9540 65156 9568
rect 65150 9528 65156 9540
rect 65225 9537 65237 9571
rect 65208 9531 65237 9537
rect 65208 9528 65214 9531
rect 64874 9500 64880 9512
rect 64800 9472 64880 9500
rect 64874 9460 64880 9472
rect 64932 9460 64938 9512
rect 64966 9460 64972 9512
rect 65024 9500 65030 9512
rect 65981 9503 66039 9509
rect 65981 9500 65993 9503
rect 65024 9472 65993 9500
rect 65024 9460 65030 9472
rect 65981 9469 65993 9472
rect 66027 9469 66039 9503
rect 65981 9463 66039 9469
rect 64984 9432 65012 9460
rect 64892 9404 65012 9432
rect 64892 9373 64920 9404
rect 65058 9392 65064 9444
rect 65116 9432 65122 9444
rect 65429 9435 65487 9441
rect 65429 9432 65441 9435
rect 65116 9404 65441 9432
rect 65116 9392 65122 9404
rect 65429 9401 65441 9404
rect 65475 9401 65487 9435
rect 65429 9395 65487 9401
rect 64877 9367 64935 9373
rect 64877 9333 64889 9367
rect 64923 9333 64935 9367
rect 64877 9327 64935 9333
rect 64966 9324 64972 9376
rect 65024 9324 65030 9376
rect 65150 9324 65156 9376
rect 65208 9364 65214 9376
rect 65337 9367 65395 9373
rect 65337 9364 65349 9367
rect 65208 9336 65349 9364
rect 65208 9324 65214 9336
rect 65337 9333 65349 9336
rect 65383 9333 65395 9367
rect 65337 9327 65395 9333
rect 63572 9274 66424 9296
rect 63572 9222 65258 9274
rect 65310 9222 65322 9274
rect 65374 9222 65386 9274
rect 65438 9222 65450 9274
rect 65502 9222 65514 9274
rect 65566 9222 66424 9274
rect 63572 9200 66424 9222
rect 64601 9163 64659 9169
rect 64601 9129 64613 9163
rect 64647 9160 64659 9163
rect 64690 9160 64696 9172
rect 64647 9132 64696 9160
rect 64647 9129 64659 9132
rect 64601 9123 64659 9129
rect 64690 9120 64696 9132
rect 64748 9120 64754 9172
rect 64969 9163 65027 9169
rect 64969 9129 64981 9163
rect 65015 9160 65027 9163
rect 65058 9160 65064 9172
rect 65015 9132 65064 9160
rect 65015 9129 65027 9132
rect 64969 9123 65027 9129
rect 65058 9120 65064 9132
rect 65116 9120 65122 9172
rect 64966 8984 64972 9036
rect 65024 9024 65030 9036
rect 65978 9024 65984 9036
rect 65024 8996 65984 9024
rect 65024 8984 65030 8996
rect 65978 8984 65984 8996
rect 66036 8984 66042 9036
rect 63494 8916 63500 8968
rect 63552 8956 63558 8968
rect 64230 8956 64236 8968
rect 63552 8928 64236 8956
rect 63552 8916 63558 8928
rect 64230 8916 64236 8928
rect 64288 8916 64294 8968
rect 65058 8916 65064 8968
rect 65116 8916 65122 8968
rect 65242 8916 65248 8968
rect 65300 8956 65306 8968
rect 65702 8956 65708 8968
rect 65300 8928 65708 8956
rect 65300 8916 65306 8928
rect 65702 8916 65708 8928
rect 65760 8916 65766 8968
rect 63572 8730 66424 8752
rect 63572 8678 64338 8730
rect 64390 8678 64402 8730
rect 64454 8678 64466 8730
rect 64518 8678 64530 8730
rect 64582 8678 64594 8730
rect 64646 8678 66424 8730
rect 63572 8656 66424 8678
rect 65242 8440 65248 8492
rect 65300 8440 65306 8492
rect 65061 8415 65119 8421
rect 65061 8381 65073 8415
rect 65107 8412 65119 8415
rect 65610 8412 65616 8424
rect 65107 8384 65616 8412
rect 65107 8381 65119 8384
rect 65061 8375 65119 8381
rect 65610 8372 65616 8384
rect 65668 8372 65674 8424
rect 65794 8372 65800 8424
rect 65852 8412 65858 8424
rect 65981 8415 66039 8421
rect 65981 8412 65993 8415
rect 65852 8384 65993 8412
rect 65852 8372 65858 8384
rect 65981 8381 65993 8384
rect 66027 8381 66039 8415
rect 65981 8375 66039 8381
rect 64969 8347 65027 8353
rect 64969 8313 64981 8347
rect 65015 8344 65027 8347
rect 65429 8347 65487 8353
rect 65429 8344 65441 8347
rect 65015 8316 65441 8344
rect 65015 8313 65027 8316
rect 64969 8307 65027 8313
rect 65429 8313 65441 8316
rect 65475 8313 65487 8347
rect 65429 8307 65487 8313
rect 64598 8236 64604 8288
rect 64656 8236 64662 8288
rect 63572 8186 66424 8208
rect 63572 8134 65258 8186
rect 65310 8134 65322 8186
rect 65374 8134 65386 8186
rect 65438 8134 65450 8186
rect 65502 8134 65514 8186
rect 65566 8134 66424 8186
rect 63572 8112 66424 8134
rect 64325 8007 64383 8013
rect 64325 7973 64337 8007
rect 64371 8004 64383 8007
rect 64598 8004 64604 8016
rect 64371 7976 64604 8004
rect 64371 7973 64383 7976
rect 64325 7967 64383 7973
rect 64598 7964 64604 7976
rect 64656 7964 64662 8016
rect 66162 8004 66168 8016
rect 65550 7976 66168 8004
rect 66162 7964 66168 7976
rect 66220 7964 66226 8016
rect 64046 7896 64052 7948
rect 64104 7896 64110 7948
rect 65794 7692 65800 7744
rect 65852 7692 65858 7744
rect 63572 7642 66424 7664
rect 63572 7590 64338 7642
rect 64390 7590 64402 7642
rect 64454 7590 64466 7642
rect 64518 7590 64530 7642
rect 64582 7590 64594 7642
rect 64646 7590 66424 7642
rect 63572 7568 66424 7590
rect 65058 7488 65064 7540
rect 65116 7528 65122 7540
rect 65245 7531 65303 7537
rect 65245 7528 65257 7531
rect 65116 7500 65257 7528
rect 65116 7488 65122 7500
rect 65245 7497 65257 7500
rect 65291 7497 65303 7531
rect 65245 7491 65303 7497
rect 64874 7460 64880 7472
rect 64708 7432 64880 7460
rect 64708 7401 64736 7432
rect 64874 7420 64880 7432
rect 64932 7420 64938 7472
rect 64693 7395 64751 7401
rect 64693 7361 64705 7395
rect 64739 7361 64751 7395
rect 64693 7355 64751 7361
rect 64785 7395 64843 7401
rect 64785 7361 64797 7395
rect 64831 7392 64843 7395
rect 65794 7392 65800 7404
rect 64831 7364 65800 7392
rect 64831 7361 64843 7364
rect 64785 7355 64843 7361
rect 65794 7352 65800 7364
rect 65852 7352 65858 7404
rect 64506 7284 64512 7336
rect 64564 7324 64570 7336
rect 64877 7327 64935 7333
rect 64877 7324 64889 7327
rect 64564 7296 64889 7324
rect 64564 7284 64570 7296
rect 64877 7293 64889 7296
rect 64923 7293 64935 7327
rect 64877 7287 64935 7293
rect 65978 7284 65984 7336
rect 66036 7284 66042 7336
rect 65429 7191 65487 7197
rect 65429 7157 65441 7191
rect 65475 7188 65487 7191
rect 65610 7188 65616 7200
rect 65475 7160 65616 7188
rect 65475 7157 65487 7160
rect 65429 7151 65487 7157
rect 65610 7148 65616 7160
rect 65668 7148 65674 7200
rect 63572 7098 66424 7120
rect 63572 7046 65258 7098
rect 65310 7046 65322 7098
rect 65374 7046 65386 7098
rect 65438 7046 65450 7098
rect 65502 7046 65514 7098
rect 65566 7046 66424 7098
rect 63572 7024 66424 7046
rect 65245 6987 65303 6993
rect 65245 6953 65257 6987
rect 65291 6984 65303 6987
rect 65610 6984 65616 6996
rect 65291 6956 65616 6984
rect 65291 6953 65303 6956
rect 65245 6947 65303 6953
rect 65610 6944 65616 6956
rect 65668 6944 65674 6996
rect 62850 6808 62856 6860
rect 62908 6848 62914 6860
rect 63586 6848 63592 6860
rect 62908 6820 63592 6848
rect 62908 6808 62914 6820
rect 63586 6808 63592 6820
rect 63644 6848 63650 6860
rect 63865 6851 63923 6857
rect 63865 6848 63877 6851
rect 63644 6820 63877 6848
rect 63644 6808 63650 6820
rect 63865 6817 63877 6820
rect 63911 6817 63923 6851
rect 63865 6811 63923 6817
rect 64506 6808 64512 6860
rect 64564 6808 64570 6860
rect 64598 6808 64604 6860
rect 64656 6848 64662 6860
rect 64693 6851 64751 6857
rect 64693 6848 64705 6851
rect 64656 6820 64705 6848
rect 64656 6808 64662 6820
rect 64693 6817 64705 6820
rect 64739 6817 64751 6851
rect 64693 6811 64751 6817
rect 65150 6808 65156 6860
rect 65208 6848 65214 6860
rect 65337 6851 65395 6857
rect 65337 6848 65349 6851
rect 65208 6820 65349 6848
rect 65208 6808 65214 6820
rect 65337 6817 65349 6820
rect 65383 6817 65395 6851
rect 65337 6811 65395 6817
rect 64141 6783 64199 6789
rect 64141 6749 64153 6783
rect 64187 6780 64199 6783
rect 64966 6780 64972 6792
rect 64187 6752 64972 6780
rect 64187 6749 64199 6752
rect 64141 6743 64199 6749
rect 64966 6740 64972 6752
rect 65024 6740 65030 6792
rect 65521 6783 65579 6789
rect 65521 6749 65533 6783
rect 65567 6780 65579 6783
rect 65610 6780 65616 6792
rect 65567 6752 65616 6780
rect 65567 6749 65579 6752
rect 65521 6743 65579 6749
rect 65610 6740 65616 6752
rect 65668 6740 65674 6792
rect 64782 6604 64788 6656
rect 64840 6644 64846 6656
rect 64877 6647 64935 6653
rect 64877 6644 64889 6647
rect 64840 6616 64889 6644
rect 64840 6604 64846 6616
rect 64877 6613 64889 6616
rect 64923 6613 64935 6647
rect 64877 6607 64935 6613
rect 63572 6554 66424 6576
rect 63572 6502 64338 6554
rect 64390 6502 64402 6554
rect 64454 6502 64466 6554
rect 64518 6502 64530 6554
rect 64582 6502 64594 6554
rect 64646 6502 66424 6554
rect 63572 6480 66424 6502
rect 64693 6443 64751 6449
rect 64693 6409 64705 6443
rect 64739 6440 64751 6443
rect 66254 6440 66260 6452
rect 64739 6412 66260 6440
rect 64739 6409 64751 6412
rect 64693 6403 64751 6409
rect 66254 6400 66260 6412
rect 66312 6400 66318 6452
rect 64138 6332 64144 6384
rect 64196 6372 64202 6384
rect 64506 6372 64512 6384
rect 64196 6344 64512 6372
rect 64196 6332 64202 6344
rect 64506 6332 64512 6344
rect 64564 6332 64570 6384
rect 64049 6307 64107 6313
rect 64049 6273 64061 6307
rect 64095 6304 64107 6307
rect 64966 6304 64972 6316
rect 64095 6276 64972 6304
rect 64095 6273 64107 6276
rect 64049 6267 64107 6273
rect 64966 6264 64972 6276
rect 65024 6304 65030 6316
rect 65245 6307 65303 6313
rect 65245 6304 65257 6307
rect 65024 6276 65257 6304
rect 65024 6264 65030 6276
rect 65245 6273 65257 6276
rect 65291 6273 65303 6307
rect 65245 6267 65303 6273
rect 63954 6196 63960 6248
rect 64012 6236 64018 6248
rect 64141 6239 64199 6245
rect 64141 6236 64153 6239
rect 64012 6208 64153 6236
rect 64012 6196 64018 6208
rect 64141 6205 64153 6208
rect 64187 6205 64199 6239
rect 64141 6199 64199 6205
rect 64506 6196 64512 6248
rect 64564 6236 64570 6248
rect 65061 6239 65119 6245
rect 65061 6236 65073 6239
rect 64564 6208 65073 6236
rect 64564 6196 64570 6208
rect 65061 6205 65073 6208
rect 65107 6205 65119 6239
rect 65061 6199 65119 6205
rect 65153 6239 65211 6245
rect 65153 6205 65165 6239
rect 65199 6236 65211 6239
rect 65978 6236 65984 6248
rect 65199 6208 65984 6236
rect 65199 6205 65211 6208
rect 65153 6199 65211 6205
rect 65978 6196 65984 6208
rect 66036 6196 66042 6248
rect 64233 6171 64291 6177
rect 64233 6137 64245 6171
rect 64279 6168 64291 6171
rect 64874 6168 64880 6180
rect 64279 6140 64880 6168
rect 64279 6137 64291 6140
rect 64233 6131 64291 6137
rect 64874 6128 64880 6140
rect 64932 6128 64938 6180
rect 64322 6060 64328 6112
rect 64380 6100 64386 6112
rect 64601 6103 64659 6109
rect 64601 6100 64613 6103
rect 64380 6072 64613 6100
rect 64380 6060 64386 6072
rect 64601 6069 64613 6072
rect 64647 6069 64659 6103
rect 64601 6063 64659 6069
rect 63572 6010 66424 6032
rect 63572 5958 65258 6010
rect 65310 5958 65322 6010
rect 65374 5958 65386 6010
rect 65438 5958 65450 6010
rect 65502 5958 65514 6010
rect 65566 5958 66424 6010
rect 63572 5936 66424 5958
rect 63586 5856 63592 5908
rect 63644 5896 63650 5908
rect 64138 5896 64144 5908
rect 63644 5868 64144 5896
rect 63644 5856 63650 5868
rect 64138 5856 64144 5868
rect 64196 5856 64202 5908
rect 64322 5856 64328 5908
rect 64380 5856 64386 5908
rect 64506 5856 64512 5908
rect 64564 5896 64570 5908
rect 64693 5899 64751 5905
rect 64693 5896 64705 5899
rect 64564 5868 64705 5896
rect 64564 5856 64570 5868
rect 64693 5865 64705 5868
rect 64739 5865 64751 5899
rect 64693 5859 64751 5865
rect 63586 5720 63592 5772
rect 63644 5760 63650 5772
rect 64233 5763 64291 5769
rect 64233 5760 64245 5763
rect 63644 5732 64245 5760
rect 63644 5720 63650 5732
rect 64233 5729 64245 5732
rect 64279 5729 64291 5763
rect 64233 5723 64291 5729
rect 64322 5652 64328 5704
rect 64380 5692 64386 5704
rect 64417 5695 64475 5701
rect 64417 5692 64429 5695
rect 64380 5664 64429 5692
rect 64380 5652 64386 5664
rect 64417 5661 64429 5664
rect 64463 5661 64475 5695
rect 64417 5655 64475 5661
rect 63865 5559 63923 5565
rect 63865 5525 63877 5559
rect 63911 5556 63923 5559
rect 63954 5556 63960 5568
rect 63911 5528 63960 5556
rect 63911 5525 63923 5528
rect 63865 5519 63923 5525
rect 63954 5516 63960 5528
rect 64012 5516 64018 5568
rect 63572 5466 66424 5488
rect 63572 5414 64338 5466
rect 64390 5414 64402 5466
rect 64454 5414 64466 5466
rect 64518 5414 64530 5466
rect 64582 5414 64594 5466
rect 64646 5414 66424 5466
rect 63572 5392 66424 5414
rect 65797 5355 65855 5361
rect 65797 5321 65809 5355
rect 65843 5352 65855 5355
rect 65978 5352 65984 5364
rect 65843 5324 65984 5352
rect 65843 5321 65855 5324
rect 65797 5315 65855 5321
rect 65978 5312 65984 5324
rect 66036 5312 66042 5364
rect 64046 5176 64052 5228
rect 64104 5176 64110 5228
rect 64325 5219 64383 5225
rect 64325 5185 64337 5219
rect 64371 5216 64383 5219
rect 64782 5216 64788 5228
rect 64371 5188 64788 5216
rect 64371 5185 64383 5188
rect 64325 5179 64383 5185
rect 64782 5176 64788 5188
rect 64840 5176 64846 5228
rect 65702 5080 65708 5092
rect 65550 5052 65708 5080
rect 65702 5040 65708 5052
rect 65760 5080 65766 5092
rect 66162 5080 66168 5092
rect 65760 5052 66168 5080
rect 65760 5040 65766 5052
rect 66162 5040 66168 5052
rect 66220 5040 66226 5092
rect 63572 4922 66424 4944
rect 63572 4870 65258 4922
rect 65310 4870 65322 4922
rect 65374 4870 65386 4922
rect 65438 4870 65450 4922
rect 65502 4870 65514 4922
rect 65566 4870 66424 4922
rect 63572 4848 66424 4870
rect 64874 4768 64880 4820
rect 64932 4808 64938 4820
rect 65150 4808 65156 4820
rect 64932 4780 65156 4808
rect 64932 4768 64938 4780
rect 65150 4768 65156 4780
rect 65208 4808 65214 4820
rect 65613 4811 65671 4817
rect 65613 4808 65625 4811
rect 65208 4780 65625 4808
rect 65208 4768 65214 4780
rect 65613 4777 65625 4780
rect 65659 4777 65671 4811
rect 65613 4771 65671 4777
rect 65702 4740 65708 4752
rect 65366 4712 65708 4740
rect 65702 4700 65708 4712
rect 65760 4700 65766 4752
rect 63862 4632 63868 4684
rect 63920 4632 63926 4684
rect 64141 4607 64199 4613
rect 64141 4573 64153 4607
rect 64187 4604 64199 4607
rect 64690 4604 64696 4616
rect 64187 4576 64696 4604
rect 64187 4573 64199 4576
rect 64141 4567 64199 4573
rect 64690 4564 64696 4576
rect 64748 4564 64754 4616
rect 63572 4378 66424 4400
rect 63572 4326 64338 4378
rect 64390 4326 64402 4378
rect 64454 4326 64466 4378
rect 64518 4326 64530 4378
rect 64582 4326 64594 4378
rect 64646 4326 66424 4378
rect 63572 4304 66424 4326
rect 63954 4224 63960 4276
rect 64012 4264 64018 4276
rect 64122 4267 64180 4273
rect 64122 4264 64134 4267
rect 64012 4236 64134 4264
rect 64012 4224 64018 4236
rect 64122 4233 64134 4236
rect 64168 4233 64180 4267
rect 64122 4227 64180 4233
rect 63865 4063 63923 4069
rect 63865 4029 63877 4063
rect 63911 4029 63923 4063
rect 63865 4023 63923 4029
rect 63880 3992 63908 4023
rect 64046 3992 64052 4004
rect 63880 3964 64052 3992
rect 64046 3952 64052 3964
rect 64104 3952 64110 4004
rect 66438 3992 66444 4004
rect 65366 3964 66444 3992
rect 66438 3952 66444 3964
rect 66496 3952 66502 4004
rect 64138 3884 64144 3936
rect 64196 3924 64202 3936
rect 65613 3927 65671 3933
rect 65613 3924 65625 3927
rect 64196 3896 65625 3924
rect 64196 3884 64202 3896
rect 65613 3893 65625 3896
rect 65659 3893 65671 3927
rect 65613 3887 65671 3893
rect 63572 3834 66424 3856
rect 63572 3782 65258 3834
rect 65310 3782 65322 3834
rect 65374 3782 65386 3834
rect 65438 3782 65450 3834
rect 65502 3782 65514 3834
rect 65566 3782 66424 3834
rect 63572 3760 66424 3782
rect 64138 3680 64144 3732
rect 64196 3680 64202 3732
rect 64601 3723 64659 3729
rect 64601 3689 64613 3723
rect 64647 3720 64659 3723
rect 65153 3723 65211 3729
rect 65153 3720 65165 3723
rect 64647 3692 65165 3720
rect 64647 3689 64659 3692
rect 64601 3683 64659 3689
rect 65153 3689 65165 3692
rect 65199 3689 65211 3723
rect 65153 3683 65211 3689
rect 63494 3612 63500 3664
rect 63552 3652 63558 3664
rect 63862 3652 63868 3664
rect 63552 3624 63868 3652
rect 63552 3612 63558 3624
rect 63862 3612 63868 3624
rect 63920 3652 63926 3664
rect 64233 3655 64291 3661
rect 64233 3652 64245 3655
rect 63920 3624 64245 3652
rect 63920 3612 63926 3624
rect 64233 3621 64245 3624
rect 64279 3621 64291 3655
rect 64233 3615 64291 3621
rect 65058 3544 65064 3596
rect 65116 3544 65122 3596
rect 64049 3519 64107 3525
rect 64049 3485 64061 3519
rect 64095 3485 64107 3519
rect 64049 3479 64107 3485
rect 65337 3519 65395 3525
rect 65337 3485 65349 3519
rect 65383 3516 65395 3519
rect 65610 3516 65616 3528
rect 65383 3488 65616 3516
rect 65383 3485 65395 3488
rect 65337 3479 65395 3485
rect 64064 3448 64092 3479
rect 65610 3476 65616 3488
rect 65668 3476 65674 3528
rect 64966 3448 64972 3460
rect 64064 3420 64972 3448
rect 64966 3408 64972 3420
rect 65024 3408 65030 3460
rect 64690 3340 64696 3392
rect 64748 3340 64754 3392
rect 63572 3290 66424 3312
rect 63572 3238 64338 3290
rect 64390 3238 64402 3290
rect 64454 3238 64466 3290
rect 64518 3238 64530 3290
rect 64582 3238 64594 3290
rect 64646 3238 66424 3290
rect 63572 3216 66424 3238
rect 63862 3136 63868 3188
rect 63920 3136 63926 3188
rect 64046 3000 64052 3052
rect 64104 3000 64110 3052
rect 64230 2864 64236 2916
rect 64288 2904 64294 2916
rect 64325 2907 64383 2913
rect 64325 2904 64337 2907
rect 64288 2876 64337 2904
rect 64288 2864 64294 2876
rect 64325 2873 64337 2876
rect 64371 2873 64383 2907
rect 65702 2904 65708 2916
rect 65550 2876 65708 2904
rect 64325 2867 64383 2873
rect 65702 2864 65708 2876
rect 65760 2864 65766 2916
rect 65794 2796 65800 2848
rect 65852 2796 65858 2848
rect 63572 2746 66424 2768
rect 63572 2694 65258 2746
rect 65310 2694 65322 2746
rect 65374 2694 65386 2746
rect 65438 2694 65450 2746
rect 65502 2694 65514 2746
rect 65566 2694 66424 2746
rect 63572 2672 66424 2694
rect 63586 2592 63592 2644
rect 63644 2632 63650 2644
rect 63865 2635 63923 2641
rect 63865 2632 63877 2635
rect 63644 2604 63877 2632
rect 63644 2592 63650 2604
rect 63865 2601 63877 2604
rect 63911 2601 63923 2635
rect 63865 2595 63923 2601
rect 64693 2635 64751 2641
rect 64693 2601 64705 2635
rect 64739 2632 64751 2635
rect 64966 2632 64972 2644
rect 64739 2604 64972 2632
rect 64739 2601 64751 2604
rect 64693 2595 64751 2601
rect 64966 2592 64972 2604
rect 65024 2592 65030 2644
rect 65153 2635 65211 2641
rect 65153 2601 65165 2635
rect 65199 2632 65211 2635
rect 66070 2632 66076 2644
rect 65199 2604 66076 2632
rect 65199 2601 65211 2604
rect 65153 2595 65211 2601
rect 66070 2592 66076 2604
rect 66128 2592 66134 2644
rect 64138 2456 64144 2508
rect 64196 2496 64202 2508
rect 64417 2499 64475 2505
rect 64417 2496 64429 2499
rect 64196 2468 64429 2496
rect 64196 2456 64202 2468
rect 64417 2465 64429 2468
rect 64463 2465 64475 2499
rect 64417 2459 64475 2465
rect 65150 2456 65156 2508
rect 65208 2496 65214 2508
rect 65245 2499 65303 2505
rect 65245 2496 65257 2499
rect 65208 2468 65257 2496
rect 65208 2456 65214 2468
rect 65245 2465 65257 2468
rect 65291 2465 65303 2499
rect 65245 2459 65303 2465
rect 64322 2388 64328 2440
rect 64380 2428 64386 2440
rect 64690 2428 64696 2440
rect 64380 2400 64696 2428
rect 64380 2388 64386 2400
rect 64690 2388 64696 2400
rect 64748 2428 64754 2440
rect 65337 2431 65395 2437
rect 64748 2400 64874 2428
rect 64748 2388 64754 2400
rect 64846 2360 64874 2400
rect 65337 2397 65349 2431
rect 65383 2397 65395 2431
rect 65337 2391 65395 2397
rect 65352 2360 65380 2391
rect 64846 2332 65380 2360
rect 64782 2252 64788 2304
rect 64840 2252 64846 2304
rect 63572 2202 66424 2224
rect 63572 2150 64338 2202
rect 64390 2150 64402 2202
rect 64454 2150 64466 2202
rect 64518 2150 64530 2202
rect 64582 2150 64594 2202
rect 64646 2150 66424 2202
rect 63572 2128 66424 2150
rect 65058 2048 65064 2100
rect 65116 2088 65122 2100
rect 65429 2091 65487 2097
rect 65429 2088 65441 2091
rect 65116 2060 65441 2088
rect 65116 2048 65122 2060
rect 65429 2057 65441 2060
rect 65475 2057 65487 2091
rect 65429 2051 65487 2057
rect 48958 1980 48964 2032
rect 49016 2020 49022 2032
rect 63034 2020 63040 2032
rect 49016 1992 63040 2020
rect 49016 1980 49022 1992
rect 63034 1980 63040 1992
rect 63092 1980 63098 2032
rect 65337 2023 65395 2029
rect 65337 1989 65349 2023
rect 65383 2020 65395 2023
rect 65886 2020 65892 2032
rect 65383 1992 65892 2020
rect 65383 1989 65395 1992
rect 65337 1983 65395 1989
rect 65886 1980 65892 1992
rect 65944 1980 65950 2032
rect 49602 1912 49608 1964
rect 49660 1952 49666 1964
rect 62482 1952 62488 1964
rect 49660 1924 62488 1952
rect 49660 1912 49666 1924
rect 62482 1912 62488 1924
rect 62540 1912 62546 1964
rect 64690 1912 64696 1964
rect 64748 1912 64754 1964
rect 64877 1955 64935 1961
rect 64877 1921 64889 1955
rect 64923 1952 64935 1955
rect 65794 1952 65800 1964
rect 64923 1924 65800 1952
rect 64923 1921 64935 1924
rect 64877 1915 64935 1921
rect 65794 1912 65800 1924
rect 65852 1912 65858 1964
rect 49694 1844 49700 1896
rect 49752 1884 49758 1896
rect 63770 1884 63776 1896
rect 49752 1856 63776 1884
rect 49752 1844 49758 1856
rect 63770 1844 63776 1856
rect 63828 1844 63834 1896
rect 65150 1844 65156 1896
rect 65208 1884 65214 1896
rect 65981 1887 66039 1893
rect 65981 1884 65993 1887
rect 65208 1856 65993 1884
rect 65208 1844 65214 1856
rect 65981 1853 65993 1856
rect 66027 1853 66039 1887
rect 65981 1847 66039 1853
rect 64690 1776 64696 1828
rect 64748 1816 64754 1828
rect 64966 1816 64972 1828
rect 64748 1788 64972 1816
rect 64748 1776 64754 1788
rect 64966 1776 64972 1788
rect 65024 1776 65030 1828
rect 63572 1658 66424 1680
rect 63572 1606 65258 1658
rect 65310 1606 65322 1658
rect 65374 1606 65386 1658
rect 65438 1606 65450 1658
rect 65502 1606 65514 1658
rect 65566 1606 66424 1658
rect 63572 1584 66424 1606
rect 64690 1504 64696 1556
rect 64748 1504 64754 1556
rect 64782 1504 64788 1556
rect 64840 1544 64846 1556
rect 65245 1547 65303 1553
rect 65245 1544 65257 1547
rect 64840 1516 65257 1544
rect 64840 1504 64846 1516
rect 65245 1513 65257 1516
rect 65291 1513 65303 1547
rect 65245 1507 65303 1513
rect 64230 1368 64236 1420
rect 64288 1408 64294 1420
rect 64288 1380 64828 1408
rect 64288 1368 64294 1380
rect 64800 1281 64828 1380
rect 65150 1368 65156 1420
rect 65208 1368 65214 1420
rect 65429 1343 65487 1349
rect 65429 1309 65441 1343
rect 65475 1340 65487 1343
rect 65610 1340 65616 1352
rect 65475 1312 65616 1340
rect 65475 1309 65487 1312
rect 65429 1303 65487 1309
rect 65610 1300 65616 1312
rect 65668 1300 65674 1352
rect 64785 1275 64843 1281
rect 64785 1241 64797 1275
rect 64831 1241 64843 1275
rect 64785 1235 64843 1241
rect 63572 1114 66424 1136
rect 63572 1062 64338 1114
rect 64390 1062 64402 1114
rect 64454 1062 64466 1114
rect 64518 1062 64530 1114
rect 64582 1062 64594 1114
rect 64646 1062 66424 1114
rect 63572 1040 66424 1062
rect 65150 960 65156 1012
rect 65208 1000 65214 1012
rect 65429 1003 65487 1009
rect 65429 1000 65441 1003
rect 65208 972 65441 1000
rect 65208 960 65214 972
rect 65429 969 65441 972
rect 65475 969 65487 1003
rect 65429 963 65487 969
rect 65794 824 65800 876
rect 65852 864 65858 876
rect 65981 867 66039 873
rect 65981 864 65993 867
rect 65852 836 65993 864
rect 65852 824 65858 836
rect 65981 833 65993 836
rect 66027 833 66039 867
rect 65981 827 66039 833
rect 63572 570 66424 592
rect 63572 518 65258 570
rect 65310 518 65322 570
rect 65374 518 65386 570
rect 65438 518 65450 570
rect 65502 518 65514 570
rect 65566 518 66424 570
rect 63572 496 66424 518
<< via1 >>
rect 21272 44956 21324 45008
rect 39396 44956 39448 45008
rect 15108 44752 15160 44804
rect 22836 44752 22888 44804
rect 14556 44684 14608 44736
rect 21456 44684 21508 44736
rect 22008 44684 22060 44736
rect 23296 44684 23348 44736
rect 26424 44684 26476 44736
rect 29092 44684 29144 44736
rect 32404 44684 32456 44736
rect 1998 44582 2050 44634
rect 2062 44582 2114 44634
rect 2126 44582 2178 44634
rect 2190 44582 2242 44634
rect 2254 44582 2306 44634
rect 49998 44582 50050 44634
rect 50062 44582 50114 44634
rect 50126 44582 50178 44634
rect 50190 44582 50242 44634
rect 50254 44582 50306 44634
rect 6184 44523 6236 44532
rect 6184 44489 6193 44523
rect 6193 44489 6227 44523
rect 6227 44489 6236 44523
rect 6184 44480 6236 44489
rect 6736 44523 6788 44532
rect 6736 44489 6745 44523
rect 6745 44489 6779 44523
rect 6779 44489 6788 44523
rect 6736 44480 6788 44489
rect 7288 44523 7340 44532
rect 7288 44489 7297 44523
rect 7297 44489 7331 44523
rect 7331 44489 7340 44523
rect 7288 44480 7340 44489
rect 7840 44523 7892 44532
rect 7840 44489 7849 44523
rect 7849 44489 7883 44523
rect 7883 44489 7892 44523
rect 7840 44480 7892 44489
rect 8392 44523 8444 44532
rect 8392 44489 8401 44523
rect 8401 44489 8435 44523
rect 8435 44489 8444 44523
rect 8392 44480 8444 44489
rect 8944 44523 8996 44532
rect 8944 44489 8953 44523
rect 8953 44489 8987 44523
rect 8987 44489 8996 44523
rect 8944 44480 8996 44489
rect 9496 44523 9548 44532
rect 9496 44489 9505 44523
rect 9505 44489 9539 44523
rect 9539 44489 9548 44523
rect 9496 44480 9548 44489
rect 10048 44523 10100 44532
rect 10048 44489 10057 44523
rect 10057 44489 10091 44523
rect 10091 44489 10100 44523
rect 10048 44480 10100 44489
rect 10508 44523 10560 44532
rect 10508 44489 10517 44523
rect 10517 44489 10551 44523
rect 10551 44489 10560 44523
rect 10508 44480 10560 44489
rect 10784 44523 10836 44532
rect 10784 44489 10793 44523
rect 10793 44489 10827 44523
rect 10827 44489 10836 44523
rect 10784 44480 10836 44489
rect 11152 44523 11204 44532
rect 11152 44489 11161 44523
rect 11161 44489 11195 44523
rect 11195 44489 11204 44523
rect 11152 44480 11204 44489
rect 11428 44523 11480 44532
rect 11428 44489 11437 44523
rect 11437 44489 11471 44523
rect 11471 44489 11480 44523
rect 11428 44480 11480 44489
rect 11704 44523 11756 44532
rect 11704 44489 11713 44523
rect 11713 44489 11747 44523
rect 11747 44489 11756 44523
rect 11704 44480 11756 44489
rect 12532 44523 12584 44532
rect 12532 44489 12541 44523
rect 12541 44489 12575 44523
rect 12575 44489 12584 44523
rect 12532 44480 12584 44489
rect 15200 44480 15252 44532
rect 18420 44480 18472 44532
rect 13820 44412 13872 44464
rect 16488 44412 16540 44464
rect 19708 44412 19760 44464
rect 17224 44344 17276 44396
rect 19524 44344 19576 44396
rect 20076 44523 20128 44532
rect 20076 44489 20085 44523
rect 20085 44489 20119 44523
rect 20119 44489 20128 44523
rect 20076 44480 20128 44489
rect 19892 44412 19944 44464
rect 21640 44412 21692 44464
rect 14372 44276 14424 44328
rect 14556 44319 14608 44328
rect 14556 44285 14565 44319
rect 14565 44285 14599 44319
rect 14599 44285 14608 44319
rect 14556 44276 14608 44285
rect 15108 44319 15160 44328
rect 15108 44285 15117 44319
rect 15117 44285 15151 44319
rect 15151 44285 15160 44319
rect 15108 44276 15160 44285
rect 15384 44319 15436 44328
rect 15384 44285 15393 44319
rect 15393 44285 15427 44319
rect 15427 44285 15436 44319
rect 15384 44276 15436 44285
rect 17776 44276 17828 44328
rect 19708 44276 19760 44328
rect 21916 44344 21968 44396
rect 22008 44344 22060 44396
rect 22560 44276 22612 44328
rect 11612 44140 11664 44192
rect 13728 44183 13780 44192
rect 13728 44149 13737 44183
rect 13737 44149 13771 44183
rect 13771 44149 13780 44183
rect 13728 44140 13780 44149
rect 14096 44208 14148 44260
rect 14740 44140 14792 44192
rect 17592 44208 17644 44260
rect 17684 44208 17736 44260
rect 20720 44208 20772 44260
rect 26332 44480 26384 44532
rect 26424 44480 26476 44532
rect 23020 44412 23072 44464
rect 24768 44344 24820 44396
rect 25044 44344 25096 44396
rect 25688 44387 25740 44396
rect 25688 44353 25697 44387
rect 25697 44353 25731 44387
rect 25731 44353 25740 44387
rect 25688 44344 25740 44353
rect 27344 44344 27396 44396
rect 28080 44344 28132 44396
rect 28724 44344 28776 44396
rect 32404 44523 32456 44532
rect 32404 44489 32413 44523
rect 32413 44489 32447 44523
rect 32447 44489 32456 44523
rect 32404 44480 32456 44489
rect 32956 44480 33008 44532
rect 27988 44319 28040 44328
rect 27988 44285 27997 44319
rect 27997 44285 28031 44319
rect 28031 44285 28040 44319
rect 27988 44276 28040 44285
rect 31024 44319 31076 44328
rect 31024 44285 31033 44319
rect 31033 44285 31067 44319
rect 31067 44285 31076 44319
rect 31024 44276 31076 44285
rect 35164 44344 35216 44396
rect 38292 44344 38344 44396
rect 15936 44183 15988 44192
rect 15936 44149 15945 44183
rect 15945 44149 15979 44183
rect 15979 44149 15988 44183
rect 15936 44140 15988 44149
rect 16856 44140 16908 44192
rect 18144 44140 18196 44192
rect 18972 44140 19024 44192
rect 19800 44140 19852 44192
rect 21180 44140 21232 44192
rect 21732 44140 21784 44192
rect 25228 44208 25280 44260
rect 25504 44208 25556 44260
rect 26884 44251 26936 44260
rect 26884 44217 26893 44251
rect 26893 44217 26927 44251
rect 26927 44217 26936 44251
rect 26884 44208 26936 44217
rect 23480 44140 23532 44192
rect 23664 44183 23716 44192
rect 23664 44149 23673 44183
rect 23673 44149 23707 44183
rect 23707 44149 23716 44183
rect 23664 44140 23716 44149
rect 24216 44140 24268 44192
rect 24676 44183 24728 44192
rect 24676 44149 24685 44183
rect 24685 44149 24719 44183
rect 24719 44149 24728 44183
rect 24676 44140 24728 44149
rect 24768 44183 24820 44192
rect 24768 44149 24777 44183
rect 24777 44149 24811 44183
rect 24811 44149 24820 44183
rect 24768 44140 24820 44149
rect 25688 44140 25740 44192
rect 26516 44140 26568 44192
rect 27896 44140 27948 44192
rect 28816 44140 28868 44192
rect 33416 44276 33468 44328
rect 34336 44276 34388 44328
rect 35256 44276 35308 44328
rect 36728 44276 36780 44328
rect 38844 44319 38896 44328
rect 38844 44285 38853 44319
rect 38853 44285 38887 44319
rect 38887 44285 38896 44319
rect 38844 44276 38896 44285
rect 31300 44140 31352 44192
rect 33324 44208 33376 44260
rect 37740 44208 37792 44260
rect 39948 44276 40000 44328
rect 40316 44276 40368 44328
rect 39304 44208 39356 44260
rect 43444 44412 43496 44464
rect 41420 44344 41472 44396
rect 41236 44276 41288 44328
rect 44364 44344 44416 44396
rect 43352 44319 43404 44328
rect 43352 44285 43361 44319
rect 43361 44285 43395 44319
rect 43395 44285 43404 44319
rect 43352 44276 43404 44285
rect 44180 44276 44232 44328
rect 47400 44412 47452 44464
rect 46112 44344 46164 44396
rect 45928 44276 45980 44328
rect 52736 44276 52788 44328
rect 33232 44183 33284 44192
rect 33232 44149 33241 44183
rect 33241 44149 33275 44183
rect 33275 44149 33284 44183
rect 33232 44140 33284 44149
rect 34428 44140 34480 44192
rect 34520 44140 34572 44192
rect 35532 44140 35584 44192
rect 35808 44183 35860 44192
rect 35808 44149 35817 44183
rect 35817 44149 35851 44183
rect 35851 44149 35860 44183
rect 35808 44140 35860 44149
rect 36544 44140 36596 44192
rect 38200 44140 38252 44192
rect 39488 44140 39540 44192
rect 40868 44140 40920 44192
rect 44732 44251 44784 44260
rect 44732 44217 44741 44251
rect 44741 44217 44775 44251
rect 44775 44217 44784 44251
rect 44732 44208 44784 44217
rect 41420 44183 41472 44192
rect 41420 44149 41429 44183
rect 41429 44149 41463 44183
rect 41463 44149 41472 44183
rect 41420 44140 41472 44149
rect 42156 44140 42208 44192
rect 42340 44183 42392 44192
rect 42340 44149 42349 44183
rect 42349 44149 42383 44183
rect 42383 44149 42392 44183
rect 42340 44140 42392 44149
rect 42524 44140 42576 44192
rect 45376 44140 45428 44192
rect 46020 44140 46072 44192
rect 46664 44140 46716 44192
rect 47400 44251 47452 44260
rect 47400 44217 47409 44251
rect 47409 44217 47443 44251
rect 47443 44217 47452 44251
rect 47400 44208 47452 44217
rect 48044 44208 48096 44260
rect 53840 44140 53892 44192
rect 2918 44038 2970 44090
rect 2982 44038 3034 44090
rect 3046 44038 3098 44090
rect 3110 44038 3162 44090
rect 3174 44038 3226 44090
rect 50918 44038 50970 44090
rect 50982 44038 51034 44090
rect 51046 44038 51098 44090
rect 51110 44038 51162 44090
rect 51174 44038 51226 44090
rect 14648 43936 14700 43988
rect 12532 43868 12584 43920
rect 12808 43843 12860 43852
rect 12808 43809 12817 43843
rect 12817 43809 12851 43843
rect 12851 43809 12860 43843
rect 12808 43800 12860 43809
rect 11612 43775 11664 43784
rect 11612 43741 11621 43775
rect 11621 43741 11655 43775
rect 11655 43741 11664 43775
rect 11612 43732 11664 43741
rect 11704 43732 11756 43784
rect 12256 43664 12308 43716
rect 13728 43868 13780 43920
rect 15200 43868 15252 43920
rect 15936 43936 15988 43988
rect 17408 43936 17460 43988
rect 17776 43979 17828 43988
rect 17776 43945 17785 43979
rect 17785 43945 17819 43979
rect 17819 43945 17828 43979
rect 17776 43936 17828 43945
rect 18328 43979 18380 43988
rect 18328 43945 18337 43979
rect 18337 43945 18371 43979
rect 18371 43945 18380 43979
rect 18328 43936 18380 43945
rect 11060 43639 11112 43648
rect 11060 43605 11069 43639
rect 11069 43605 11103 43639
rect 11103 43605 11112 43639
rect 11060 43596 11112 43605
rect 12624 43596 12676 43648
rect 13820 43664 13872 43716
rect 16212 43843 16264 43852
rect 16212 43809 16221 43843
rect 16221 43809 16255 43843
rect 16255 43809 16264 43843
rect 16212 43800 16264 43809
rect 14924 43732 14976 43784
rect 13636 43639 13688 43648
rect 13636 43605 13645 43639
rect 13645 43605 13679 43639
rect 13679 43605 13688 43639
rect 13636 43596 13688 43605
rect 14464 43639 14516 43648
rect 14464 43605 14473 43639
rect 14473 43605 14507 43639
rect 14507 43605 14516 43639
rect 14464 43596 14516 43605
rect 15936 43596 15988 43648
rect 17132 43596 17184 43648
rect 19340 43868 19392 43920
rect 20720 43936 20772 43988
rect 21548 43936 21600 43988
rect 21732 43979 21784 43988
rect 21732 43945 21741 43979
rect 21741 43945 21775 43979
rect 21775 43945 21784 43979
rect 21732 43936 21784 43945
rect 24676 43936 24728 43988
rect 24952 43936 25004 43988
rect 19432 43800 19484 43852
rect 21640 43843 21692 43852
rect 21640 43809 21649 43843
rect 21649 43809 21683 43843
rect 21683 43809 21692 43843
rect 21640 43800 21692 43809
rect 21916 43868 21968 43920
rect 23020 43868 23072 43920
rect 23664 43868 23716 43920
rect 24860 43868 24912 43920
rect 32956 43936 33008 43988
rect 33416 43979 33468 43988
rect 33416 43945 33425 43979
rect 33425 43945 33459 43979
rect 33459 43945 33468 43979
rect 33416 43936 33468 43945
rect 36544 43979 36596 43988
rect 36544 43945 36553 43979
rect 36553 43945 36587 43979
rect 36587 43945 36596 43979
rect 36544 43936 36596 43945
rect 36728 43979 36780 43988
rect 36728 43945 36737 43979
rect 36737 43945 36771 43979
rect 36771 43945 36780 43979
rect 36728 43936 36780 43945
rect 27896 43868 27948 43920
rect 29092 43868 29144 43920
rect 22284 43800 22336 43852
rect 26240 43800 26292 43852
rect 26884 43800 26936 43852
rect 30564 43800 30616 43852
rect 32220 43868 32272 43920
rect 33324 43868 33376 43920
rect 35256 43868 35308 43920
rect 36360 43868 36412 43920
rect 37740 43868 37792 43920
rect 38200 43911 38252 43920
rect 38200 43877 38209 43911
rect 38209 43877 38243 43911
rect 38243 43877 38252 43911
rect 38200 43868 38252 43877
rect 35440 43843 35492 43852
rect 35440 43809 35449 43843
rect 35449 43809 35483 43843
rect 35483 43809 35492 43843
rect 35440 43800 35492 43809
rect 39396 43936 39448 43988
rect 41236 43936 41288 43988
rect 44732 43936 44784 43988
rect 17592 43732 17644 43784
rect 17868 43775 17920 43784
rect 17868 43741 17877 43775
rect 17877 43741 17911 43775
rect 17911 43741 17920 43775
rect 17868 43732 17920 43741
rect 21088 43775 21140 43784
rect 21088 43741 21097 43775
rect 21097 43741 21131 43775
rect 21131 43741 21140 43775
rect 21088 43732 21140 43741
rect 22100 43732 22152 43784
rect 22376 43775 22428 43784
rect 22376 43741 22385 43775
rect 22385 43741 22419 43775
rect 22419 43741 22428 43775
rect 22376 43732 22428 43741
rect 22744 43732 22796 43784
rect 23388 43775 23440 43784
rect 23388 43741 23397 43775
rect 23397 43741 23431 43775
rect 23431 43741 23440 43775
rect 23388 43732 23440 43741
rect 18420 43596 18472 43648
rect 19432 43596 19484 43648
rect 19708 43596 19760 43648
rect 21456 43707 21508 43716
rect 21456 43673 21465 43707
rect 21465 43673 21499 43707
rect 21499 43673 21508 43707
rect 21456 43664 21508 43673
rect 21824 43664 21876 43716
rect 26792 43732 26844 43784
rect 27252 43732 27304 43784
rect 26608 43664 26660 43716
rect 29552 43732 29604 43784
rect 29920 43732 29972 43784
rect 33232 43732 33284 43784
rect 20076 43596 20128 43648
rect 20168 43596 20220 43648
rect 21088 43596 21140 43648
rect 22468 43596 22520 43648
rect 25872 43596 25924 43648
rect 26056 43639 26108 43648
rect 26056 43605 26065 43639
rect 26065 43605 26099 43639
rect 26099 43605 26108 43639
rect 26056 43596 26108 43605
rect 31024 43596 31076 43648
rect 31760 43596 31812 43648
rect 34152 43732 34204 43784
rect 35348 43732 35400 43784
rect 35808 43732 35860 43784
rect 38476 43775 38528 43784
rect 38476 43741 38485 43775
rect 38485 43741 38519 43775
rect 38519 43741 38528 43775
rect 38476 43732 38528 43741
rect 40960 43775 41012 43784
rect 40960 43741 40969 43775
rect 40969 43741 41003 43775
rect 41003 43741 41012 43775
rect 40960 43732 41012 43741
rect 41236 43775 41288 43784
rect 41236 43741 41245 43775
rect 41245 43741 41279 43775
rect 41279 43741 41288 43775
rect 41236 43732 41288 43741
rect 42156 43911 42208 43920
rect 42156 43877 42165 43911
rect 42165 43877 42199 43911
rect 42199 43877 42208 43911
rect 42156 43868 42208 43877
rect 43444 43868 43496 43920
rect 46664 43868 46716 43920
rect 41880 43775 41932 43784
rect 41880 43741 41889 43775
rect 41889 43741 41923 43775
rect 41923 43741 41932 43775
rect 41880 43732 41932 43741
rect 43168 43732 43220 43784
rect 43904 43800 43956 43852
rect 52552 43843 52604 43852
rect 52552 43809 52561 43843
rect 52561 43809 52595 43843
rect 52595 43809 52604 43843
rect 52552 43800 52604 43809
rect 52736 43843 52788 43852
rect 52736 43809 52745 43843
rect 52745 43809 52779 43843
rect 52779 43809 52788 43843
rect 52736 43800 52788 43809
rect 44916 43732 44968 43784
rect 47400 43732 47452 43784
rect 47492 43775 47544 43784
rect 47492 43741 47501 43775
rect 47501 43741 47535 43775
rect 47535 43741 47544 43775
rect 47492 43732 47544 43741
rect 47952 43732 48004 43784
rect 44180 43664 44232 43716
rect 44456 43664 44508 43716
rect 66352 43800 66404 43852
rect 35072 43596 35124 43648
rect 35256 43639 35308 43648
rect 35256 43605 35265 43639
rect 35265 43605 35299 43639
rect 35299 43605 35308 43639
rect 35256 43596 35308 43605
rect 35532 43639 35584 43648
rect 35532 43605 35541 43639
rect 35541 43605 35575 43639
rect 35575 43605 35584 43639
rect 35532 43596 35584 43605
rect 38568 43639 38620 43648
rect 38568 43605 38577 43639
rect 38577 43605 38611 43639
rect 38611 43605 38620 43639
rect 38568 43596 38620 43605
rect 43812 43639 43864 43648
rect 43812 43605 43821 43639
rect 43821 43605 43855 43639
rect 43855 43605 43864 43639
rect 43812 43596 43864 43605
rect 47308 43596 47360 43648
rect 48228 43596 48280 43648
rect 51908 43596 51960 43648
rect 53196 43596 53248 43648
rect 1998 43494 2050 43546
rect 2062 43494 2114 43546
rect 2126 43494 2178 43546
rect 2190 43494 2242 43546
rect 2254 43494 2306 43546
rect 49998 43494 50050 43546
rect 50062 43494 50114 43546
rect 50126 43494 50178 43546
rect 50190 43494 50242 43546
rect 50254 43494 50306 43546
rect 15384 43392 15436 43444
rect 17500 43435 17552 43444
rect 17500 43401 17509 43435
rect 17509 43401 17543 43435
rect 17543 43401 17552 43435
rect 17500 43392 17552 43401
rect 19524 43392 19576 43444
rect 20536 43392 20588 43444
rect 18052 43324 18104 43376
rect 20076 43324 20128 43376
rect 22560 43435 22612 43444
rect 22560 43401 22569 43435
rect 22569 43401 22603 43435
rect 22603 43401 22612 43435
rect 22560 43392 22612 43401
rect 23388 43392 23440 43444
rect 25780 43392 25832 43444
rect 28816 43435 28868 43444
rect 28816 43401 28825 43435
rect 28825 43401 28859 43435
rect 28859 43401 28868 43435
rect 28816 43392 28868 43401
rect 28908 43392 28960 43444
rect 23296 43324 23348 43376
rect 25228 43324 25280 43376
rect 26424 43324 26476 43376
rect 13636 43256 13688 43308
rect 10692 43231 10744 43240
rect 10692 43197 10701 43231
rect 10701 43197 10735 43231
rect 10735 43197 10744 43231
rect 10692 43188 10744 43197
rect 11244 43120 11296 43172
rect 15384 43231 15436 43240
rect 15384 43197 15393 43231
rect 15393 43197 15427 43231
rect 15427 43197 15436 43231
rect 15384 43188 15436 43197
rect 18144 43231 18196 43240
rect 18144 43197 18153 43231
rect 18153 43197 18187 43231
rect 18187 43197 18196 43231
rect 18144 43188 18196 43197
rect 18420 43299 18472 43308
rect 18420 43265 18429 43299
rect 18429 43265 18463 43299
rect 18463 43265 18472 43299
rect 18420 43256 18472 43265
rect 13820 43120 13872 43172
rect 15936 43163 15988 43172
rect 15936 43129 15945 43163
rect 15945 43129 15979 43163
rect 15979 43129 15988 43163
rect 15936 43120 15988 43129
rect 17684 43120 17736 43172
rect 18972 43163 19024 43172
rect 18972 43129 18981 43163
rect 18981 43129 19015 43163
rect 19015 43129 19024 43163
rect 18972 43120 19024 43129
rect 20352 43120 20404 43172
rect 12716 43052 12768 43104
rect 12992 43052 13044 43104
rect 13728 43052 13780 43104
rect 15568 43052 15620 43104
rect 17776 43095 17828 43104
rect 17776 43061 17785 43095
rect 17785 43061 17819 43095
rect 17819 43061 17828 43095
rect 17776 43052 17828 43061
rect 19984 43052 20036 43104
rect 26240 43256 26292 43308
rect 27436 43324 27488 43376
rect 28080 43324 28132 43376
rect 29552 43435 29604 43444
rect 29552 43401 29561 43435
rect 29561 43401 29595 43435
rect 29595 43401 29604 43435
rect 29552 43392 29604 43401
rect 23480 43188 23532 43240
rect 23664 43231 23716 43240
rect 23664 43197 23673 43231
rect 23673 43197 23707 43231
rect 23707 43197 23716 43231
rect 23664 43188 23716 43197
rect 26056 43188 26108 43240
rect 28540 43256 28592 43308
rect 29920 43324 29972 43376
rect 34152 43435 34204 43444
rect 34152 43401 34161 43435
rect 34161 43401 34195 43435
rect 34195 43401 34204 43435
rect 34152 43392 34204 43401
rect 34428 43392 34480 43444
rect 36360 43435 36412 43444
rect 36360 43401 36369 43435
rect 36369 43401 36403 43435
rect 36403 43401 36412 43435
rect 36360 43392 36412 43401
rect 40960 43392 41012 43444
rect 42340 43392 42392 43444
rect 43812 43392 43864 43444
rect 28356 43231 28408 43240
rect 28356 43197 28365 43231
rect 28365 43197 28399 43231
rect 28399 43197 28408 43231
rect 28356 43188 28408 43197
rect 29920 43231 29972 43240
rect 29920 43197 29929 43231
rect 29929 43197 29963 43231
rect 29963 43197 29972 43231
rect 29920 43188 29972 43197
rect 21180 43120 21232 43172
rect 21640 43120 21692 43172
rect 24216 43120 24268 43172
rect 24860 43120 24912 43172
rect 22008 43052 22060 43104
rect 22836 43095 22888 43104
rect 22836 43061 22845 43095
rect 22845 43061 22879 43095
rect 22879 43061 22888 43095
rect 22836 43052 22888 43061
rect 23020 43095 23072 43104
rect 23020 43061 23029 43095
rect 23029 43061 23063 43095
rect 23063 43061 23072 43095
rect 23020 43052 23072 43061
rect 25412 43052 25464 43104
rect 25872 43052 25924 43104
rect 27528 43163 27580 43172
rect 27528 43129 27537 43163
rect 27537 43129 27571 43163
rect 27571 43129 27580 43163
rect 27528 43120 27580 43129
rect 28908 43120 28960 43172
rect 30288 43188 30340 43240
rect 31760 43299 31812 43308
rect 31760 43265 31769 43299
rect 31769 43265 31803 43299
rect 31803 43265 31812 43299
rect 31760 43256 31812 43265
rect 35440 43324 35492 43376
rect 39396 43324 39448 43376
rect 33324 43256 33376 43308
rect 26240 43052 26292 43104
rect 27344 43095 27396 43104
rect 27344 43061 27353 43095
rect 27353 43061 27387 43095
rect 27387 43061 27396 43095
rect 27344 43052 27396 43061
rect 27436 43052 27488 43104
rect 31208 43120 31260 43172
rect 30012 43095 30064 43104
rect 30012 43061 30021 43095
rect 30021 43061 30055 43095
rect 30055 43061 30064 43095
rect 30012 43052 30064 43061
rect 30564 43095 30616 43104
rect 30564 43061 30573 43095
rect 30573 43061 30607 43095
rect 30607 43061 30616 43095
rect 30564 43052 30616 43061
rect 31300 43052 31352 43104
rect 35164 43256 35216 43308
rect 34520 43231 34572 43240
rect 34520 43197 34529 43231
rect 34529 43197 34563 43231
rect 34563 43197 34572 43231
rect 34520 43188 34572 43197
rect 35256 43188 35308 43240
rect 32036 43163 32088 43172
rect 32036 43129 32045 43163
rect 32045 43129 32079 43163
rect 32079 43129 32088 43163
rect 32036 43120 32088 43129
rect 32496 43120 32548 43172
rect 34428 43120 34480 43172
rect 34796 43052 34848 43104
rect 35348 43052 35400 43104
rect 38292 43256 38344 43308
rect 40132 43256 40184 43308
rect 41236 43324 41288 43376
rect 37740 43120 37792 43172
rect 37924 43120 37976 43172
rect 38568 43231 38620 43240
rect 38568 43197 38577 43231
rect 38577 43197 38611 43231
rect 38611 43197 38620 43231
rect 38568 43188 38620 43197
rect 40316 43231 40368 43240
rect 40316 43197 40325 43231
rect 40325 43197 40359 43231
rect 40359 43197 40368 43231
rect 40316 43188 40368 43197
rect 41420 43299 41472 43308
rect 41420 43265 41429 43299
rect 41429 43265 41463 43299
rect 41463 43265 41472 43299
rect 41420 43256 41472 43265
rect 43352 43324 43404 43376
rect 47492 43392 47544 43444
rect 49516 43392 49568 43444
rect 52552 43392 52604 43444
rect 38844 43120 38896 43172
rect 39396 43163 39448 43172
rect 39396 43129 39405 43163
rect 39405 43129 39439 43163
rect 39439 43129 39448 43163
rect 39396 43120 39448 43129
rect 43076 43188 43128 43240
rect 43996 43299 44048 43308
rect 43996 43265 44005 43299
rect 44005 43265 44039 43299
rect 44039 43265 44048 43299
rect 43996 43256 44048 43265
rect 44088 43299 44140 43308
rect 44088 43265 44097 43299
rect 44097 43265 44131 43299
rect 44131 43265 44140 43299
rect 44088 43256 44140 43265
rect 45376 43299 45428 43308
rect 45376 43265 45385 43299
rect 45385 43265 45419 43299
rect 45419 43265 45428 43299
rect 45376 43256 45428 43265
rect 45928 43256 45980 43308
rect 46848 43299 46900 43308
rect 46848 43265 46857 43299
rect 46857 43265 46891 43299
rect 46891 43265 46900 43299
rect 46848 43256 46900 43265
rect 47308 43299 47360 43308
rect 47308 43265 47317 43299
rect 47317 43265 47351 43299
rect 47351 43265 47360 43299
rect 47308 43256 47360 43265
rect 51264 43256 51316 43308
rect 52552 43256 52604 43308
rect 44824 43188 44876 43240
rect 46940 43188 46992 43240
rect 53840 43231 53892 43240
rect 53840 43197 53849 43231
rect 53849 43197 53883 43231
rect 53883 43197 53892 43231
rect 53840 43188 53892 43197
rect 38384 43052 38436 43104
rect 39304 43052 39356 43104
rect 39580 43052 39632 43104
rect 40408 43095 40460 43104
rect 40408 43061 40417 43095
rect 40417 43061 40451 43095
rect 40451 43061 40460 43095
rect 40408 43052 40460 43061
rect 41788 43052 41840 43104
rect 41972 43163 42024 43172
rect 41972 43129 41981 43163
rect 41981 43129 42015 43163
rect 42015 43129 42024 43163
rect 41972 43120 42024 43129
rect 46664 43120 46716 43172
rect 48964 43120 49016 43172
rect 53196 43120 53248 43172
rect 51540 43052 51592 43104
rect 52460 43095 52512 43104
rect 52460 43061 52469 43095
rect 52469 43061 52503 43095
rect 52503 43061 52512 43095
rect 52460 43052 52512 43061
rect 53380 43095 53432 43104
rect 53380 43061 53389 43095
rect 53389 43061 53423 43095
rect 53423 43061 53432 43095
rect 53380 43052 53432 43061
rect 60648 43052 60700 43104
rect 2918 42950 2970 43002
rect 2982 42950 3034 43002
rect 3046 42950 3098 43002
rect 3110 42950 3162 43002
rect 3174 42950 3226 43002
rect 50918 42950 50970 43002
rect 50982 42950 51034 43002
rect 51046 42950 51098 43002
rect 51110 42950 51162 43002
rect 51174 42950 51226 43002
rect 11244 42848 11296 42900
rect 11704 42891 11756 42900
rect 11704 42857 11713 42891
rect 11713 42857 11747 42891
rect 11747 42857 11756 42891
rect 11704 42848 11756 42857
rect 14648 42848 14700 42900
rect 15200 42891 15252 42900
rect 15200 42857 15209 42891
rect 15209 42857 15243 42891
rect 15243 42857 15252 42891
rect 15200 42848 15252 42857
rect 16856 42891 16908 42900
rect 16856 42857 16865 42891
rect 16865 42857 16899 42891
rect 16899 42857 16908 42891
rect 16856 42848 16908 42857
rect 17684 42848 17736 42900
rect 13820 42780 13872 42832
rect 15568 42823 15620 42832
rect 15568 42789 15577 42823
rect 15577 42789 15611 42823
rect 15611 42789 15620 42823
rect 15568 42780 15620 42789
rect 12716 42712 12768 42764
rect 15844 42712 15896 42764
rect 16488 42780 16540 42832
rect 17132 42780 17184 42832
rect 17776 42780 17828 42832
rect 19340 42891 19392 42900
rect 19340 42857 19349 42891
rect 19349 42857 19383 42891
rect 19383 42857 19392 42891
rect 19340 42848 19392 42857
rect 19984 42848 20036 42900
rect 20444 42891 20496 42900
rect 20444 42857 20453 42891
rect 20453 42857 20487 42891
rect 20487 42857 20496 42891
rect 20444 42848 20496 42857
rect 20536 42891 20588 42900
rect 20536 42857 20545 42891
rect 20545 42857 20579 42891
rect 20579 42857 20588 42891
rect 20536 42848 20588 42857
rect 9496 42687 9548 42696
rect 9496 42653 9505 42687
rect 9505 42653 9539 42687
rect 9539 42653 9548 42687
rect 9496 42644 9548 42653
rect 12624 42644 12676 42696
rect 12808 42687 12860 42696
rect 12808 42653 12817 42687
rect 12817 42653 12851 42687
rect 12851 42653 12860 42687
rect 12808 42644 12860 42653
rect 14464 42644 14516 42696
rect 8944 42551 8996 42560
rect 8944 42517 8953 42551
rect 8953 42517 8987 42551
rect 8987 42517 8996 42551
rect 8944 42508 8996 42517
rect 13176 42508 13228 42560
rect 13544 42508 13596 42560
rect 16672 42644 16724 42696
rect 16948 42687 17000 42696
rect 16948 42653 16957 42687
rect 16957 42653 16991 42687
rect 16991 42653 17000 42687
rect 16948 42644 17000 42653
rect 17132 42687 17184 42696
rect 17132 42653 17141 42687
rect 17141 42653 17175 42687
rect 17175 42653 17184 42687
rect 17132 42644 17184 42653
rect 17316 42755 17368 42764
rect 17316 42721 17325 42755
rect 17325 42721 17359 42755
rect 17359 42721 17368 42755
rect 17316 42712 17368 42721
rect 17592 42755 17644 42764
rect 17592 42721 17601 42755
rect 17601 42721 17635 42755
rect 17635 42721 17644 42755
rect 17592 42712 17644 42721
rect 22652 42780 22704 42832
rect 22836 42780 22888 42832
rect 23480 42848 23532 42900
rect 24952 42848 25004 42900
rect 25780 42891 25832 42900
rect 25780 42857 25789 42891
rect 25789 42857 25823 42891
rect 25823 42857 25832 42891
rect 25780 42848 25832 42857
rect 25964 42848 26016 42900
rect 26240 42891 26292 42900
rect 26240 42857 26249 42891
rect 26249 42857 26283 42891
rect 26283 42857 26292 42891
rect 26240 42848 26292 42857
rect 26332 42848 26384 42900
rect 27344 42848 27396 42900
rect 27988 42891 28040 42900
rect 27988 42857 27997 42891
rect 27997 42857 28031 42891
rect 28031 42857 28040 42891
rect 27988 42848 28040 42857
rect 30012 42848 30064 42900
rect 30564 42848 30616 42900
rect 31760 42848 31812 42900
rect 32496 42848 32548 42900
rect 32588 42848 32640 42900
rect 33048 42891 33100 42900
rect 33048 42857 33057 42891
rect 33057 42857 33091 42891
rect 33091 42857 33100 42891
rect 33048 42848 33100 42857
rect 34336 42891 34388 42900
rect 34336 42857 34345 42891
rect 34345 42857 34379 42891
rect 34379 42857 34388 42891
rect 34336 42848 34388 42857
rect 34796 42891 34848 42900
rect 34796 42857 34805 42891
rect 34805 42857 34839 42891
rect 34839 42857 34848 42891
rect 34796 42848 34848 42857
rect 36728 42848 36780 42900
rect 39488 42891 39540 42900
rect 39488 42857 39497 42891
rect 39497 42857 39531 42891
rect 39531 42857 39540 42891
rect 39488 42848 39540 42857
rect 24860 42780 24912 42832
rect 20352 42712 20404 42764
rect 22560 42712 22612 42764
rect 25044 42755 25096 42764
rect 16028 42576 16080 42628
rect 20536 42644 20588 42696
rect 21364 42687 21416 42696
rect 21364 42653 21373 42687
rect 21373 42653 21407 42687
rect 21407 42653 21416 42687
rect 21364 42644 21416 42653
rect 25044 42721 25053 42755
rect 25053 42721 25087 42755
rect 25087 42721 25096 42755
rect 25044 42712 25096 42721
rect 16304 42551 16356 42560
rect 16304 42517 16313 42551
rect 16313 42517 16347 42551
rect 16347 42517 16356 42551
rect 16304 42508 16356 42517
rect 16396 42508 16448 42560
rect 21272 42576 21324 42628
rect 22192 42576 22244 42628
rect 24676 42644 24728 42696
rect 17592 42508 17644 42560
rect 20168 42508 20220 42560
rect 20536 42508 20588 42560
rect 22376 42508 22428 42560
rect 22560 42508 22612 42560
rect 22836 42508 22888 42560
rect 24952 42576 25004 42628
rect 24216 42508 24268 42560
rect 25136 42687 25188 42696
rect 25136 42653 25145 42687
rect 25145 42653 25179 42687
rect 25179 42653 25188 42687
rect 25136 42644 25188 42653
rect 25228 42644 25280 42696
rect 26056 42712 26108 42764
rect 25688 42687 25740 42696
rect 25688 42653 25697 42687
rect 25697 42653 25731 42687
rect 25731 42653 25740 42687
rect 26516 42712 26568 42764
rect 30656 42780 30708 42832
rect 36176 42823 36228 42832
rect 36176 42789 36185 42823
rect 36185 42789 36219 42823
rect 36219 42789 36228 42823
rect 36176 42780 36228 42789
rect 36360 42780 36412 42832
rect 27528 42712 27580 42764
rect 28540 42712 28592 42764
rect 25688 42644 25740 42653
rect 28080 42687 28132 42696
rect 28080 42653 28089 42687
rect 28089 42653 28123 42687
rect 28123 42653 28132 42687
rect 28080 42644 28132 42653
rect 28448 42644 28500 42696
rect 29460 42644 29512 42696
rect 31024 42712 31076 42764
rect 31300 42712 31352 42764
rect 30472 42687 30524 42696
rect 30472 42653 30481 42687
rect 30481 42653 30515 42687
rect 30515 42653 30524 42687
rect 30472 42644 30524 42653
rect 31852 42644 31904 42696
rect 32312 42712 32364 42764
rect 33232 42644 33284 42696
rect 33508 42755 33560 42764
rect 33508 42721 33517 42755
rect 33517 42721 33551 42755
rect 33551 42721 33560 42755
rect 33508 42712 33560 42721
rect 34060 42712 34112 42764
rect 36636 42712 36688 42764
rect 38108 42712 38160 42764
rect 33600 42687 33652 42696
rect 33600 42653 33609 42687
rect 33609 42653 33643 42687
rect 33643 42653 33652 42687
rect 33600 42644 33652 42653
rect 26516 42576 26568 42628
rect 26700 42551 26752 42560
rect 26700 42517 26709 42551
rect 26709 42517 26743 42551
rect 26743 42517 26752 42551
rect 26700 42508 26752 42517
rect 26884 42508 26936 42560
rect 32036 42576 32088 42628
rect 33416 42576 33468 42628
rect 34980 42644 35032 42696
rect 35532 42644 35584 42696
rect 36820 42687 36872 42696
rect 35348 42576 35400 42628
rect 36820 42653 36829 42687
rect 36829 42653 36863 42687
rect 36863 42653 36872 42687
rect 36820 42644 36872 42653
rect 37188 42644 37240 42696
rect 38384 42644 38436 42696
rect 38752 42644 38804 42696
rect 40408 42848 40460 42900
rect 41144 42848 41196 42900
rect 41972 42848 42024 42900
rect 42524 42848 42576 42900
rect 43996 42848 44048 42900
rect 46020 42848 46072 42900
rect 46756 42891 46808 42900
rect 46756 42857 46765 42891
rect 46765 42857 46799 42891
rect 46799 42857 46808 42891
rect 46756 42848 46808 42857
rect 47400 42848 47452 42900
rect 48228 42891 48280 42900
rect 48228 42857 48237 42891
rect 48237 42857 48271 42891
rect 48271 42857 48280 42891
rect 48228 42848 48280 42857
rect 51540 42848 51592 42900
rect 52460 42848 52512 42900
rect 40592 42687 40644 42696
rect 40592 42653 40601 42687
rect 40601 42653 40635 42687
rect 40635 42653 40644 42687
rect 40592 42644 40644 42653
rect 40776 42687 40828 42696
rect 40776 42653 40785 42687
rect 40785 42653 40819 42687
rect 40819 42653 40828 42687
rect 40776 42644 40828 42653
rect 43168 42780 43220 42832
rect 46664 42780 46716 42832
rect 46848 42780 46900 42832
rect 54024 42780 54076 42832
rect 41420 42712 41472 42764
rect 41788 42712 41840 42764
rect 44088 42712 44140 42764
rect 37832 42576 37884 42628
rect 38476 42576 38528 42628
rect 41420 42576 41472 42628
rect 36452 42508 36504 42560
rect 37464 42551 37516 42560
rect 37464 42517 37473 42551
rect 37473 42517 37507 42551
rect 37507 42517 37516 42551
rect 37464 42508 37516 42517
rect 38200 42551 38252 42560
rect 38200 42517 38209 42551
rect 38209 42517 38243 42551
rect 38243 42517 38252 42551
rect 38200 42508 38252 42517
rect 38844 42508 38896 42560
rect 40040 42508 40092 42560
rect 40592 42508 40644 42560
rect 41880 42687 41932 42696
rect 41880 42653 41889 42687
rect 41889 42653 41923 42687
rect 41923 42653 41932 42687
rect 41880 42644 41932 42653
rect 42156 42687 42208 42696
rect 42156 42653 42165 42687
rect 42165 42653 42199 42687
rect 42199 42653 42208 42687
rect 42156 42644 42208 42653
rect 42524 42644 42576 42696
rect 44180 42687 44232 42696
rect 44180 42653 44189 42687
rect 44189 42653 44223 42687
rect 44223 42653 44232 42687
rect 44180 42644 44232 42653
rect 47400 42755 47452 42764
rect 47400 42721 47409 42755
rect 47409 42721 47443 42755
rect 47443 42721 47452 42755
rect 47400 42712 47452 42721
rect 44916 42644 44968 42696
rect 45284 42687 45336 42696
rect 45284 42653 45293 42687
rect 45293 42653 45327 42687
rect 45327 42653 45336 42687
rect 45284 42644 45336 42653
rect 46848 42644 46900 42696
rect 46296 42576 46348 42628
rect 48412 42687 48464 42696
rect 48412 42653 48421 42687
rect 48421 42653 48455 42687
rect 48455 42653 48464 42687
rect 48412 42644 48464 42653
rect 43260 42508 43312 42560
rect 43628 42551 43680 42560
rect 43628 42517 43637 42551
rect 43637 42517 43671 42551
rect 43671 42517 43680 42551
rect 43628 42508 43680 42517
rect 46756 42508 46808 42560
rect 51724 42687 51776 42696
rect 51724 42653 51733 42687
rect 51733 42653 51767 42687
rect 51767 42653 51776 42687
rect 51724 42644 51776 42653
rect 51908 42687 51960 42696
rect 51908 42653 51917 42687
rect 51917 42653 51951 42687
rect 51951 42653 51960 42687
rect 51908 42644 51960 42653
rect 51540 42576 51592 42628
rect 52460 42687 52512 42696
rect 52460 42653 52469 42687
rect 52469 42653 52503 42687
rect 52503 42653 52512 42687
rect 52460 42644 52512 42653
rect 52828 42644 52880 42696
rect 51908 42508 51960 42560
rect 52920 42508 52972 42560
rect 1998 42406 2050 42458
rect 2062 42406 2114 42458
rect 2126 42406 2178 42458
rect 2190 42406 2242 42458
rect 2254 42406 2306 42458
rect 49998 42406 50050 42458
rect 50062 42406 50114 42458
rect 50126 42406 50178 42458
rect 50190 42406 50242 42458
rect 50254 42406 50306 42458
rect 11704 42347 11756 42356
rect 11704 42313 11713 42347
rect 11713 42313 11747 42347
rect 11747 42313 11756 42347
rect 11704 42304 11756 42313
rect 12532 42347 12584 42356
rect 12532 42313 12541 42347
rect 12541 42313 12575 42347
rect 12575 42313 12584 42347
rect 12532 42304 12584 42313
rect 15384 42304 15436 42356
rect 16028 42304 16080 42356
rect 16304 42304 16356 42356
rect 8392 42168 8444 42220
rect 11520 42168 11572 42220
rect 12992 42211 13044 42220
rect 12992 42177 13001 42211
rect 13001 42177 13035 42211
rect 13035 42177 13044 42211
rect 12992 42168 13044 42177
rect 13176 42211 13228 42220
rect 13176 42177 13185 42211
rect 13185 42177 13219 42211
rect 13219 42177 13228 42211
rect 13176 42168 13228 42177
rect 16948 42304 17000 42356
rect 17868 42304 17920 42356
rect 17960 42236 18012 42288
rect 16396 42168 16448 42220
rect 16672 42168 16724 42220
rect 9680 42143 9732 42152
rect 9680 42109 9689 42143
rect 9689 42109 9723 42143
rect 9723 42109 9732 42143
rect 9680 42100 9732 42109
rect 13728 42143 13780 42152
rect 13728 42109 13737 42143
rect 13737 42109 13771 42143
rect 13771 42109 13780 42143
rect 13728 42100 13780 42109
rect 8576 41964 8628 42016
rect 11060 41964 11112 42016
rect 12256 42032 12308 42084
rect 12716 42032 12768 42084
rect 13636 42032 13688 42084
rect 17684 42100 17736 42152
rect 18052 42211 18104 42220
rect 18052 42177 18061 42211
rect 18061 42177 18095 42211
rect 18095 42177 18104 42211
rect 18052 42168 18104 42177
rect 19800 42347 19852 42356
rect 19800 42313 19809 42347
rect 19809 42313 19843 42347
rect 19843 42313 19852 42347
rect 19800 42304 19852 42313
rect 20444 42304 20496 42356
rect 24768 42347 24820 42356
rect 24768 42313 24777 42347
rect 24777 42313 24811 42347
rect 24811 42313 24820 42347
rect 24768 42304 24820 42313
rect 24952 42304 25004 42356
rect 22284 42236 22336 42288
rect 20536 42168 20588 42220
rect 22008 42211 22060 42220
rect 22008 42177 22017 42211
rect 22017 42177 22051 42211
rect 22051 42177 22060 42211
rect 22008 42168 22060 42177
rect 22560 42211 22612 42220
rect 22560 42177 22569 42211
rect 22569 42177 22603 42211
rect 22603 42177 22612 42211
rect 22560 42168 22612 42177
rect 25228 42236 25280 42288
rect 25964 42304 26016 42356
rect 28356 42347 28408 42356
rect 28356 42313 28365 42347
rect 28365 42313 28399 42347
rect 28399 42313 28408 42347
rect 28356 42304 28408 42313
rect 33048 42304 33100 42356
rect 33232 42347 33284 42356
rect 33232 42313 33241 42347
rect 33241 42313 33275 42347
rect 33275 42313 33284 42347
rect 33232 42304 33284 42313
rect 33508 42304 33560 42356
rect 36176 42304 36228 42356
rect 36452 42304 36504 42356
rect 18328 42100 18380 42152
rect 19340 42100 19392 42152
rect 22100 42100 22152 42152
rect 12440 41964 12492 42016
rect 14372 42007 14424 42016
rect 14372 41973 14381 42007
rect 14381 41973 14415 42007
rect 14415 41973 14424 42007
rect 14372 41964 14424 41973
rect 15476 41964 15528 42016
rect 17960 42075 18012 42084
rect 17960 42041 17969 42075
rect 17969 42041 18003 42075
rect 18003 42041 18012 42075
rect 17960 42032 18012 42041
rect 20444 42032 20496 42084
rect 21456 42032 21508 42084
rect 21824 42032 21876 42084
rect 24032 42168 24084 42220
rect 28080 42236 28132 42288
rect 28816 42236 28868 42288
rect 23020 42100 23072 42152
rect 23756 42100 23808 42152
rect 26608 42211 26660 42220
rect 26608 42177 26617 42211
rect 26617 42177 26651 42211
rect 26651 42177 26660 42211
rect 26608 42168 26660 42177
rect 27436 42168 27488 42220
rect 32128 42168 32180 42220
rect 32220 42168 32272 42220
rect 33232 42168 33284 42220
rect 35348 42236 35400 42288
rect 34428 42168 34480 42220
rect 37464 42168 37516 42220
rect 38384 42211 38436 42220
rect 38384 42177 38393 42211
rect 38393 42177 38427 42211
rect 38427 42177 38436 42211
rect 38384 42168 38436 42177
rect 40316 42168 40368 42220
rect 40776 42304 40828 42356
rect 43904 42304 43956 42356
rect 44272 42304 44324 42356
rect 45284 42304 45336 42356
rect 49700 42304 49752 42356
rect 45928 42236 45980 42288
rect 44088 42168 44140 42220
rect 45836 42168 45888 42220
rect 46756 42168 46808 42220
rect 47768 42168 47820 42220
rect 49148 42168 49200 42220
rect 51632 42304 51684 42356
rect 51724 42304 51776 42356
rect 52460 42304 52512 42356
rect 53196 42304 53248 42356
rect 59268 42304 59320 42356
rect 51724 42168 51776 42220
rect 52644 42211 52696 42220
rect 52644 42177 52653 42211
rect 52653 42177 52687 42211
rect 52687 42177 52696 42211
rect 52644 42168 52696 42177
rect 53380 42236 53432 42288
rect 62672 42236 62724 42288
rect 53932 42168 53984 42220
rect 25044 42100 25096 42152
rect 28448 42100 28500 42152
rect 29092 42100 29144 42152
rect 31760 42100 31812 42152
rect 35072 42143 35124 42152
rect 35072 42109 35081 42143
rect 35081 42109 35115 42143
rect 35115 42109 35124 42143
rect 35072 42100 35124 42109
rect 35624 42100 35676 42152
rect 37740 42143 37792 42152
rect 37740 42109 37749 42143
rect 37749 42109 37783 42143
rect 37783 42109 37792 42143
rect 37740 42100 37792 42109
rect 38200 42143 38252 42152
rect 38200 42109 38209 42143
rect 38209 42109 38243 42143
rect 38243 42109 38252 42143
rect 38200 42100 38252 42109
rect 41420 42100 41472 42152
rect 44456 42100 44508 42152
rect 45100 42100 45152 42152
rect 52368 42100 52420 42152
rect 52552 42100 52604 42152
rect 53380 42143 53432 42152
rect 53380 42109 53389 42143
rect 53389 42109 53423 42143
rect 53423 42109 53432 42143
rect 53380 42100 53432 42109
rect 53840 42100 53892 42152
rect 63040 42100 63092 42152
rect 17040 41964 17092 42016
rect 17224 41964 17276 42016
rect 17592 41964 17644 42016
rect 17868 41964 17920 42016
rect 19708 41964 19760 42016
rect 22284 41964 22336 42016
rect 22744 41964 22796 42016
rect 23296 41964 23348 42016
rect 25412 41964 25464 42016
rect 26884 42075 26936 42084
rect 26884 42041 26893 42075
rect 26893 42041 26927 42075
rect 26927 42041 26936 42075
rect 26884 42032 26936 42041
rect 25780 41964 25832 42016
rect 28264 41964 28316 42016
rect 32864 42032 32916 42084
rect 35900 42032 35952 42084
rect 36084 42032 36136 42084
rect 30380 41964 30432 42016
rect 31852 41964 31904 42016
rect 33232 41964 33284 42016
rect 33784 41964 33836 42016
rect 37188 41964 37240 42016
rect 39580 42075 39632 42084
rect 39580 42041 39589 42075
rect 39589 42041 39623 42075
rect 39623 42041 39632 42075
rect 39580 42032 39632 42041
rect 40960 42032 41012 42084
rect 41512 42075 41564 42084
rect 41512 42041 41521 42075
rect 41521 42041 41555 42075
rect 41555 42041 41564 42075
rect 41512 42032 41564 42041
rect 41880 42075 41932 42084
rect 41880 42041 41889 42075
rect 41889 42041 41923 42075
rect 41923 42041 41932 42075
rect 41880 42032 41932 42041
rect 43168 42032 43220 42084
rect 41144 41964 41196 42016
rect 43444 42032 43496 42084
rect 44272 42032 44324 42084
rect 46296 42032 46348 42084
rect 45836 41964 45888 42016
rect 46020 42007 46072 42016
rect 46020 41973 46029 42007
rect 46029 41973 46063 42007
rect 46063 41973 46072 42007
rect 46020 41964 46072 41973
rect 48044 42032 48096 42084
rect 48320 42032 48372 42084
rect 49884 42032 49936 42084
rect 51356 42032 51408 42084
rect 53196 42032 53248 42084
rect 54024 42075 54076 42084
rect 54024 42041 54033 42075
rect 54033 42041 54067 42075
rect 54067 42041 54076 42075
rect 54024 42032 54076 42041
rect 55772 42075 55824 42084
rect 55772 42041 55781 42075
rect 55781 42041 55815 42075
rect 55815 42041 55824 42075
rect 55772 42032 55824 42041
rect 48136 41964 48188 42016
rect 48504 41964 48556 42016
rect 49792 41964 49844 42016
rect 50436 42007 50488 42016
rect 50436 41973 50445 42007
rect 50445 41973 50479 42007
rect 50479 41973 50488 42007
rect 50436 41964 50488 41973
rect 50712 41964 50764 42016
rect 52460 41964 52512 42016
rect 52644 41964 52696 42016
rect 56324 41964 56376 42016
rect 2918 41862 2970 41914
rect 2982 41862 3034 41914
rect 3046 41862 3098 41914
rect 3110 41862 3162 41914
rect 3174 41862 3226 41914
rect 50918 41862 50970 41914
rect 50982 41862 51034 41914
rect 51046 41862 51098 41914
rect 51110 41862 51162 41914
rect 51174 41862 51226 41914
rect 9496 41803 9548 41812
rect 9496 41769 9505 41803
rect 9505 41769 9539 41803
rect 9539 41769 9548 41803
rect 9496 41760 9548 41769
rect 14372 41760 14424 41812
rect 18420 41760 18472 41812
rect 18788 41760 18840 41812
rect 8300 41692 8352 41744
rect 10324 41692 10376 41744
rect 13820 41692 13872 41744
rect 16764 41692 16816 41744
rect 17040 41735 17092 41744
rect 17040 41701 17049 41735
rect 17049 41701 17083 41735
rect 17083 41701 17092 41735
rect 17040 41692 17092 41701
rect 17224 41692 17276 41744
rect 20168 41735 20220 41744
rect 20168 41701 20177 41735
rect 20177 41701 20211 41735
rect 20211 41701 20220 41735
rect 20168 41692 20220 41701
rect 22468 41803 22520 41812
rect 22468 41769 22477 41803
rect 22477 41769 22511 41803
rect 22511 41769 22520 41803
rect 22468 41760 22520 41769
rect 23664 41760 23716 41812
rect 9588 41624 9640 41676
rect 10784 41624 10836 41676
rect 8024 41599 8076 41608
rect 8024 41565 8033 41599
rect 8033 41565 8067 41599
rect 8067 41565 8076 41599
rect 8024 41556 8076 41565
rect 10232 41599 10284 41608
rect 10232 41565 10241 41599
rect 10241 41565 10275 41599
rect 10275 41565 10284 41599
rect 10232 41556 10284 41565
rect 11520 41599 11572 41608
rect 11520 41565 11529 41599
rect 11529 41565 11563 41599
rect 11563 41565 11572 41599
rect 11520 41556 11572 41565
rect 11796 41599 11848 41608
rect 11796 41565 11805 41599
rect 11805 41565 11839 41599
rect 11839 41565 11848 41599
rect 11796 41556 11848 41565
rect 12992 41556 13044 41608
rect 15568 41556 15620 41608
rect 15660 41556 15712 41608
rect 16488 41556 16540 41608
rect 16856 41599 16908 41608
rect 16856 41565 16865 41599
rect 16865 41565 16899 41599
rect 16899 41565 16908 41599
rect 16856 41556 16908 41565
rect 17132 41667 17184 41676
rect 17132 41633 17141 41667
rect 17141 41633 17175 41667
rect 17175 41633 17184 41667
rect 17132 41624 17184 41633
rect 17960 41624 18012 41676
rect 19340 41624 19392 41676
rect 23296 41735 23348 41744
rect 23296 41701 23305 41735
rect 23305 41701 23339 41735
rect 23339 41701 23348 41735
rect 23296 41692 23348 41701
rect 25136 41760 25188 41812
rect 27436 41760 27488 41812
rect 27620 41760 27672 41812
rect 26700 41735 26752 41744
rect 26700 41701 26709 41735
rect 26709 41701 26743 41735
rect 26743 41701 26752 41735
rect 26700 41692 26752 41701
rect 29460 41760 29512 41812
rect 28264 41692 28316 41744
rect 28724 41692 28776 41744
rect 33140 41760 33192 41812
rect 33232 41803 33284 41812
rect 33232 41769 33241 41803
rect 33241 41769 33275 41803
rect 33275 41769 33284 41803
rect 33232 41760 33284 41769
rect 33600 41760 33652 41812
rect 34244 41760 34296 41812
rect 36176 41760 36228 41812
rect 37188 41803 37240 41812
rect 37188 41769 37197 41803
rect 37197 41769 37231 41803
rect 37231 41769 37240 41803
rect 37188 41760 37240 41769
rect 39120 41760 39172 41812
rect 42156 41760 42208 41812
rect 42524 41760 42576 41812
rect 43352 41760 43404 41812
rect 43536 41803 43588 41812
rect 43536 41769 43545 41803
rect 43545 41769 43579 41803
rect 43579 41769 43588 41803
rect 43536 41760 43588 41769
rect 43812 41760 43864 41812
rect 43904 41760 43956 41812
rect 45008 41760 45060 41812
rect 46020 41760 46072 41812
rect 47400 41760 47452 41812
rect 29644 41692 29696 41744
rect 32036 41692 32088 41744
rect 32220 41692 32272 41744
rect 34888 41692 34940 41744
rect 18328 41599 18380 41608
rect 18328 41565 18337 41599
rect 18337 41565 18371 41599
rect 18371 41565 18380 41599
rect 18328 41556 18380 41565
rect 18420 41556 18472 41608
rect 9036 41488 9088 41540
rect 19064 41488 19116 41540
rect 22100 41556 22152 41608
rect 24860 41624 24912 41676
rect 26240 41624 26292 41676
rect 26424 41667 26476 41676
rect 26424 41633 26433 41667
rect 26433 41633 26467 41667
rect 26467 41633 26476 41667
rect 26424 41624 26476 41633
rect 29184 41624 29236 41676
rect 32864 41624 32916 41676
rect 32956 41624 33008 41676
rect 34152 41624 34204 41676
rect 22376 41556 22428 41608
rect 22560 41556 22612 41608
rect 22008 41488 22060 41540
rect 24032 41556 24084 41608
rect 25688 41556 25740 41608
rect 25964 41556 26016 41608
rect 12440 41420 12492 41472
rect 15384 41420 15436 41472
rect 17500 41463 17552 41472
rect 17500 41429 17509 41463
rect 17509 41429 17543 41463
rect 17543 41429 17552 41463
rect 17500 41420 17552 41429
rect 17960 41420 18012 41472
rect 21272 41420 21324 41472
rect 21456 41420 21508 41472
rect 22376 41420 22428 41472
rect 23296 41420 23348 41472
rect 24860 41420 24912 41472
rect 27344 41420 27396 41472
rect 28724 41599 28776 41608
rect 28724 41565 28733 41599
rect 28733 41565 28767 41599
rect 28767 41565 28776 41599
rect 28724 41556 28776 41565
rect 28816 41599 28868 41608
rect 28816 41565 28825 41599
rect 28825 41565 28859 41599
rect 28859 41565 28868 41599
rect 28816 41556 28868 41565
rect 29828 41556 29880 41608
rect 31760 41556 31812 41608
rect 32588 41556 32640 41608
rect 32680 41556 32732 41608
rect 33048 41599 33100 41608
rect 33048 41565 33057 41599
rect 33057 41565 33091 41599
rect 33091 41565 33100 41599
rect 33048 41556 33100 41565
rect 33140 41556 33192 41608
rect 34060 41599 34112 41608
rect 34060 41565 34069 41599
rect 34069 41565 34103 41599
rect 34103 41565 34112 41599
rect 34060 41556 34112 41565
rect 35992 41556 36044 41608
rect 38384 41692 38436 41744
rect 38844 41735 38896 41744
rect 38844 41701 38853 41735
rect 38853 41701 38887 41735
rect 38887 41701 38896 41735
rect 38844 41692 38896 41701
rect 40316 41692 40368 41744
rect 40500 41735 40552 41744
rect 40500 41701 40509 41735
rect 40509 41701 40543 41735
rect 40543 41701 40552 41735
rect 40500 41692 40552 41701
rect 36728 41624 36780 41676
rect 38476 41624 38528 41676
rect 39948 41624 40000 41676
rect 40960 41624 41012 41676
rect 36452 41556 36504 41608
rect 28264 41531 28316 41540
rect 28264 41497 28273 41531
rect 28273 41497 28307 41531
rect 28307 41497 28316 41531
rect 28264 41488 28316 41497
rect 28356 41488 28408 41540
rect 36544 41488 36596 41540
rect 36820 41556 36872 41608
rect 37372 41556 37424 41608
rect 30380 41420 30432 41472
rect 35808 41463 35860 41472
rect 35808 41429 35817 41463
rect 35817 41429 35851 41463
rect 35851 41429 35860 41463
rect 35808 41420 35860 41429
rect 35992 41420 36044 41472
rect 36636 41420 36688 41472
rect 38936 41420 38988 41472
rect 40224 41556 40276 41608
rect 41788 41556 41840 41608
rect 42524 41599 42576 41608
rect 42524 41565 42533 41599
rect 42533 41565 42567 41599
rect 42567 41565 42576 41599
rect 42524 41556 42576 41565
rect 40776 41488 40828 41540
rect 43168 41556 43220 41608
rect 43628 41692 43680 41744
rect 43812 41624 43864 41676
rect 44732 41624 44784 41676
rect 45928 41692 45980 41744
rect 46756 41692 46808 41744
rect 48136 41803 48188 41812
rect 48136 41769 48145 41803
rect 48145 41769 48179 41803
rect 48179 41769 48188 41803
rect 48136 41760 48188 41769
rect 48504 41803 48556 41812
rect 48504 41769 48513 41803
rect 48513 41769 48547 41803
rect 48547 41769 48556 41803
rect 48504 41760 48556 41769
rect 50436 41760 50488 41812
rect 52368 41760 52420 41812
rect 47860 41624 47912 41676
rect 40684 41420 40736 41472
rect 42708 41463 42760 41472
rect 42708 41429 42717 41463
rect 42717 41429 42751 41463
rect 42751 41429 42760 41463
rect 42708 41420 42760 41429
rect 43260 41420 43312 41472
rect 43812 41420 43864 41472
rect 44088 41420 44140 41472
rect 45836 41556 45888 41608
rect 45744 41488 45796 41540
rect 45928 41488 45980 41540
rect 46848 41556 46900 41608
rect 47584 41556 47636 41608
rect 50344 41692 50396 41744
rect 48412 41556 48464 41608
rect 49148 41556 49200 41608
rect 46940 41488 46992 41540
rect 48136 41488 48188 41540
rect 50712 41556 50764 41608
rect 52368 41556 52420 41608
rect 52920 41556 52972 41608
rect 51356 41488 51408 41540
rect 53840 41556 53892 41608
rect 55312 41599 55364 41608
rect 55312 41565 55321 41599
rect 55321 41565 55355 41599
rect 55355 41565 55364 41599
rect 55312 41556 55364 41565
rect 56508 41556 56560 41608
rect 52460 41420 52512 41472
rect 52552 41420 52604 41472
rect 52828 41420 52880 41472
rect 52920 41420 52972 41472
rect 57428 41488 57480 41540
rect 55036 41420 55088 41472
rect 1998 41318 2050 41370
rect 2062 41318 2114 41370
rect 2126 41318 2178 41370
rect 2190 41318 2242 41370
rect 2254 41318 2306 41370
rect 49998 41318 50050 41370
rect 50062 41318 50114 41370
rect 50126 41318 50178 41370
rect 50190 41318 50242 41370
rect 50254 41318 50306 41370
rect 9680 41216 9732 41268
rect 8300 41080 8352 41132
rect 8392 41123 8444 41132
rect 8392 41089 8401 41123
rect 8401 41089 8435 41123
rect 8435 41089 8444 41123
rect 8392 41080 8444 41089
rect 11796 41259 11848 41268
rect 11796 41225 11805 41259
rect 11805 41225 11839 41259
rect 11839 41225 11848 41259
rect 11796 41216 11848 41225
rect 12072 41216 12124 41268
rect 13268 41216 13320 41268
rect 15844 41216 15896 41268
rect 16488 41216 16540 41268
rect 16764 41259 16816 41268
rect 16764 41225 16773 41259
rect 16773 41225 16807 41259
rect 16807 41225 16816 41259
rect 16764 41216 16816 41225
rect 17132 41216 17184 41268
rect 17868 41216 17920 41268
rect 10232 41148 10284 41200
rect 12624 41148 12676 41200
rect 13728 41148 13780 41200
rect 11612 41080 11664 41132
rect 12900 41080 12952 41132
rect 13268 41080 13320 41132
rect 16856 41148 16908 41200
rect 17592 41148 17644 41200
rect 18604 41080 18656 41132
rect 12440 41012 12492 41064
rect 12992 41055 13044 41064
rect 12992 41021 13001 41055
rect 13001 41021 13035 41055
rect 13035 41021 13044 41055
rect 12992 41012 13044 41021
rect 8576 40944 8628 40996
rect 7748 40919 7800 40928
rect 7748 40885 7757 40919
rect 7757 40885 7791 40919
rect 7791 40885 7800 40919
rect 7748 40876 7800 40885
rect 10324 40944 10376 40996
rect 10232 40919 10284 40928
rect 10232 40885 10241 40919
rect 10241 40885 10275 40919
rect 10275 40885 10284 40919
rect 10232 40876 10284 40885
rect 11336 40876 11388 40928
rect 12440 40876 12492 40928
rect 13820 41012 13872 41064
rect 15016 41055 15068 41064
rect 15016 41021 15025 41055
rect 15025 41021 15059 41055
rect 15059 41021 15068 41055
rect 15016 41012 15068 41021
rect 18788 41080 18840 41132
rect 20168 41191 20220 41200
rect 20168 41157 20177 41191
rect 20177 41157 20211 41191
rect 20211 41157 20220 41191
rect 20168 41148 20220 41157
rect 19064 41055 19116 41064
rect 19064 41021 19073 41055
rect 19073 41021 19107 41055
rect 19107 41021 19116 41055
rect 19064 41012 19116 41021
rect 14004 40987 14056 40996
rect 14004 40953 14013 40987
rect 14013 40953 14047 40987
rect 14047 40953 14056 40987
rect 14004 40944 14056 40953
rect 15200 40944 15252 40996
rect 15752 40944 15804 40996
rect 17500 40944 17552 40996
rect 19524 40944 19576 40996
rect 23296 41148 23348 41200
rect 23756 41148 23808 41200
rect 13912 40919 13964 40928
rect 13912 40885 13921 40919
rect 13921 40885 13955 40919
rect 13955 40885 13964 40919
rect 13912 40876 13964 40885
rect 14556 40876 14608 40928
rect 17132 40876 17184 40928
rect 17408 40919 17460 40928
rect 17408 40885 17417 40919
rect 17417 40885 17451 40919
rect 17451 40885 17460 40919
rect 17408 40876 17460 40885
rect 18696 40919 18748 40928
rect 18696 40885 18705 40919
rect 18705 40885 18739 40919
rect 18739 40885 18748 40919
rect 18696 40876 18748 40885
rect 20168 40876 20220 40928
rect 22008 40987 22060 40996
rect 22008 40953 22017 40987
rect 22017 40953 22051 40987
rect 22051 40953 22060 40987
rect 22008 40944 22060 40953
rect 23020 40944 23072 40996
rect 26792 41148 26844 41200
rect 27988 41216 28040 41268
rect 30380 41216 30432 41268
rect 32956 41259 33008 41268
rect 32956 41225 32965 41259
rect 32965 41225 32999 41259
rect 32999 41225 33008 41259
rect 32956 41216 33008 41225
rect 34796 41216 34848 41268
rect 36912 41216 36964 41268
rect 43444 41216 43496 41268
rect 24492 41123 24544 41132
rect 24492 41089 24501 41123
rect 24501 41089 24535 41123
rect 24535 41089 24544 41123
rect 24492 41080 24544 41089
rect 26608 41123 26660 41132
rect 26608 41089 26617 41123
rect 26617 41089 26651 41123
rect 26651 41089 26660 41123
rect 26608 41080 26660 41089
rect 28908 41080 28960 41132
rect 30012 41080 30064 41132
rect 28356 41012 28408 41064
rect 30932 41080 30984 41132
rect 34704 41148 34756 41200
rect 36636 41191 36688 41200
rect 36636 41157 36645 41191
rect 36645 41157 36679 41191
rect 36679 41157 36688 41191
rect 36636 41148 36688 41157
rect 33232 41080 33284 41132
rect 33416 41080 33468 41132
rect 34152 41080 34204 41132
rect 35624 41080 35676 41132
rect 36728 41123 36780 41132
rect 36728 41089 36737 41123
rect 36737 41089 36771 41123
rect 36771 41089 36780 41123
rect 36728 41080 36780 41089
rect 38108 41080 38160 41132
rect 39580 41080 39632 41132
rect 40040 41148 40092 41200
rect 44088 41148 44140 41200
rect 44732 41148 44784 41200
rect 48504 41148 48556 41200
rect 49516 41148 49568 41200
rect 40132 41080 40184 41132
rect 40500 41080 40552 41132
rect 41696 41080 41748 41132
rect 30564 41012 30616 41064
rect 31484 41012 31536 41064
rect 24676 40987 24728 40996
rect 24676 40953 24685 40987
rect 24685 40953 24719 40987
rect 24719 40953 24728 40987
rect 24676 40944 24728 40953
rect 24768 40944 24820 40996
rect 32772 40944 32824 40996
rect 33692 41012 33744 41064
rect 36176 41012 36228 41064
rect 37648 41012 37700 41064
rect 38476 41012 38528 41064
rect 42248 41055 42300 41064
rect 42248 41021 42257 41055
rect 42257 41021 42291 41055
rect 42291 41021 42300 41055
rect 42248 41012 42300 41021
rect 45008 41080 45060 41132
rect 45744 41080 45796 41132
rect 46020 41123 46072 41132
rect 46020 41089 46029 41123
rect 46029 41089 46063 41123
rect 46063 41089 46072 41123
rect 46020 41080 46072 41089
rect 46296 41080 46348 41132
rect 50896 41080 50948 41132
rect 51356 41259 51408 41268
rect 51356 41225 51365 41259
rect 51365 41225 51399 41259
rect 51399 41225 51408 41259
rect 51356 41216 51408 41225
rect 53104 41216 53156 41268
rect 54024 41216 54076 41268
rect 56508 41259 56560 41268
rect 56508 41225 56517 41259
rect 56517 41225 56551 41259
rect 56551 41225 56560 41259
rect 56508 41216 56560 41225
rect 58072 41148 58124 41200
rect 66444 41148 66496 41200
rect 44272 41012 44324 41064
rect 46940 41055 46992 41064
rect 46940 41021 46949 41055
rect 46949 41021 46983 41055
rect 46983 41021 46992 41055
rect 46940 41012 46992 41021
rect 48320 41012 48372 41064
rect 49608 41055 49660 41064
rect 49608 41021 49617 41055
rect 49617 41021 49651 41055
rect 49651 41021 49660 41055
rect 49608 41012 49660 41021
rect 52644 41080 52696 41132
rect 53932 41080 53984 41132
rect 54116 41080 54168 41132
rect 64880 41080 64932 41132
rect 54760 41055 54812 41064
rect 54760 41021 54769 41055
rect 54769 41021 54803 41055
rect 54803 41021 54812 41055
rect 54760 41012 54812 41021
rect 56692 41012 56744 41064
rect 33784 40944 33836 40996
rect 22192 40876 22244 40928
rect 23756 40876 23808 40928
rect 25136 40876 25188 40928
rect 26240 40876 26292 40928
rect 29460 40919 29512 40928
rect 29460 40885 29469 40919
rect 29469 40885 29503 40919
rect 29503 40885 29512 40919
rect 29460 40876 29512 40885
rect 29920 40876 29972 40928
rect 30012 40876 30064 40928
rect 30472 40876 30524 40928
rect 31024 40876 31076 40928
rect 31392 40876 31444 40928
rect 32956 40876 33008 40928
rect 33048 40876 33100 40928
rect 33600 40919 33652 40928
rect 33600 40885 33609 40919
rect 33609 40885 33643 40919
rect 33643 40885 33652 40919
rect 33600 40876 33652 40885
rect 33968 40876 34020 40928
rect 35808 40876 35860 40928
rect 37004 40876 37056 40928
rect 37832 40876 37884 40928
rect 38108 40919 38160 40928
rect 38108 40885 38117 40919
rect 38117 40885 38151 40919
rect 38151 40885 38160 40919
rect 38108 40876 38160 40885
rect 39212 40876 39264 40928
rect 39488 40876 39540 40928
rect 39672 40919 39724 40928
rect 39672 40885 39681 40919
rect 39681 40885 39715 40919
rect 39715 40885 39724 40919
rect 39672 40876 39724 40885
rect 40500 40987 40552 40996
rect 40500 40953 40509 40987
rect 40509 40953 40543 40987
rect 40543 40953 40552 40987
rect 40500 40944 40552 40953
rect 42616 40944 42668 40996
rect 42800 40944 42852 40996
rect 43168 40944 43220 40996
rect 46020 40944 46072 40996
rect 47216 40987 47268 40996
rect 47216 40953 47225 40987
rect 47225 40953 47259 40987
rect 47259 40953 47268 40987
rect 47216 40944 47268 40953
rect 49792 40944 49844 40996
rect 41052 40876 41104 40928
rect 45100 40876 45152 40928
rect 45744 40919 45796 40928
rect 45744 40885 45753 40919
rect 45753 40885 45787 40919
rect 45787 40885 45796 40919
rect 45744 40876 45796 40885
rect 45836 40919 45888 40928
rect 45836 40885 45845 40919
rect 45845 40885 45879 40919
rect 45879 40885 45888 40919
rect 45836 40876 45888 40885
rect 48228 40876 48280 40928
rect 48688 40919 48740 40928
rect 48688 40885 48697 40919
rect 48697 40885 48731 40919
rect 48731 40885 48740 40919
rect 48688 40876 48740 40885
rect 48964 40876 49016 40928
rect 50344 40944 50396 40996
rect 52184 40944 52236 40996
rect 55036 40987 55088 40996
rect 55036 40953 55045 40987
rect 55045 40953 55079 40987
rect 55079 40953 55088 40987
rect 55036 40944 55088 40953
rect 55128 40944 55180 40996
rect 56600 40987 56652 40996
rect 56600 40953 56609 40987
rect 56609 40953 56643 40987
rect 56643 40953 56652 40987
rect 56600 40944 56652 40953
rect 57428 41055 57480 41064
rect 57428 41021 57437 41055
rect 57437 41021 57471 41055
rect 57471 41021 57480 41055
rect 57428 41012 57480 41021
rect 53472 40876 53524 40928
rect 53656 40919 53708 40928
rect 53656 40885 53665 40919
rect 53665 40885 53699 40919
rect 53699 40885 53708 40919
rect 53656 40876 53708 40885
rect 53932 40876 53984 40928
rect 54116 40876 54168 40928
rect 54668 40876 54720 40928
rect 2918 40774 2970 40826
rect 2982 40774 3034 40826
rect 3046 40774 3098 40826
rect 3110 40774 3162 40826
rect 3174 40774 3226 40826
rect 50918 40774 50970 40826
rect 50982 40774 51034 40826
rect 51046 40774 51098 40826
rect 51110 40774 51162 40826
rect 51174 40774 51226 40826
rect 8024 40672 8076 40724
rect 8944 40672 8996 40724
rect 11336 40715 11388 40724
rect 11336 40681 11345 40715
rect 11345 40681 11379 40715
rect 11379 40681 11388 40715
rect 11336 40672 11388 40681
rect 14004 40672 14056 40724
rect 15200 40715 15252 40724
rect 15200 40681 15209 40715
rect 15209 40681 15243 40715
rect 15243 40681 15252 40715
rect 15200 40672 15252 40681
rect 15476 40672 15528 40724
rect 17408 40672 17460 40724
rect 17776 40672 17828 40724
rect 9036 40647 9088 40656
rect 9036 40613 9045 40647
rect 9045 40613 9079 40647
rect 9079 40613 9088 40647
rect 9036 40604 9088 40613
rect 10324 40604 10376 40656
rect 10968 40604 11020 40656
rect 12440 40647 12492 40656
rect 12440 40613 12449 40647
rect 12449 40613 12483 40647
rect 12483 40613 12492 40647
rect 12440 40604 12492 40613
rect 12532 40604 12584 40656
rect 15016 40604 15068 40656
rect 8300 40536 8352 40588
rect 10784 40579 10836 40588
rect 10784 40545 10793 40579
rect 10793 40545 10827 40579
rect 10827 40545 10836 40579
rect 10784 40536 10836 40545
rect 11704 40536 11756 40588
rect 14556 40579 14608 40588
rect 14556 40545 14565 40579
rect 14565 40545 14599 40579
rect 14599 40545 14608 40579
rect 14556 40536 14608 40545
rect 8576 40511 8628 40520
rect 8576 40477 8585 40511
rect 8585 40477 8619 40511
rect 8619 40477 8628 40511
rect 8576 40468 8628 40477
rect 8760 40511 8812 40520
rect 8760 40477 8769 40511
rect 8769 40477 8803 40511
rect 8803 40477 8812 40511
rect 8760 40468 8812 40477
rect 10416 40468 10468 40520
rect 11244 40468 11296 40520
rect 12072 40468 12124 40520
rect 10692 40400 10744 40452
rect 13820 40468 13872 40520
rect 13912 40468 13964 40520
rect 15844 40536 15896 40588
rect 16856 40604 16908 40656
rect 18512 40579 18564 40588
rect 18512 40545 18521 40579
rect 18521 40545 18555 40579
rect 18555 40545 18564 40579
rect 18512 40536 18564 40545
rect 19248 40536 19300 40588
rect 21824 40604 21876 40656
rect 22008 40715 22060 40724
rect 22008 40681 22017 40715
rect 22017 40681 22051 40715
rect 22051 40681 22060 40715
rect 22008 40672 22060 40681
rect 23020 40672 23072 40724
rect 22652 40536 22704 40588
rect 15292 40468 15344 40520
rect 15660 40468 15712 40520
rect 15936 40468 15988 40520
rect 16488 40468 16540 40520
rect 18788 40511 18840 40520
rect 18788 40477 18797 40511
rect 18797 40477 18831 40511
rect 18831 40477 18840 40511
rect 18788 40468 18840 40477
rect 20720 40511 20772 40520
rect 20720 40477 20729 40511
rect 20729 40477 20763 40511
rect 20763 40477 20772 40511
rect 20720 40468 20772 40477
rect 17408 40400 17460 40452
rect 18328 40400 18380 40452
rect 21456 40511 21508 40520
rect 21456 40477 21465 40511
rect 21465 40477 21499 40511
rect 21499 40477 21508 40511
rect 21456 40468 21508 40477
rect 21548 40511 21600 40520
rect 21548 40477 21557 40511
rect 21557 40477 21591 40511
rect 21591 40477 21600 40511
rect 21548 40468 21600 40477
rect 21732 40468 21784 40520
rect 23204 40647 23256 40656
rect 23204 40613 23213 40647
rect 23213 40613 23247 40647
rect 23247 40613 23256 40647
rect 23204 40604 23256 40613
rect 26240 40672 26292 40724
rect 26516 40672 26568 40724
rect 23756 40647 23808 40656
rect 23756 40613 23765 40647
rect 23765 40613 23799 40647
rect 23799 40613 23808 40647
rect 23756 40604 23808 40613
rect 24768 40468 24820 40520
rect 24952 40468 25004 40520
rect 27252 40604 27304 40656
rect 27436 40672 27488 40724
rect 28264 40672 28316 40724
rect 29000 40536 29052 40588
rect 26056 40468 26108 40520
rect 27068 40511 27120 40520
rect 27068 40477 27077 40511
rect 27077 40477 27111 40511
rect 27111 40477 27120 40511
rect 27068 40468 27120 40477
rect 29920 40715 29972 40724
rect 29920 40681 29929 40715
rect 29929 40681 29963 40715
rect 29963 40681 29972 40715
rect 29920 40672 29972 40681
rect 31024 40715 31076 40724
rect 31024 40681 31033 40715
rect 31033 40681 31067 40715
rect 31067 40681 31076 40715
rect 31024 40672 31076 40681
rect 32220 40672 32272 40724
rect 32772 40672 32824 40724
rect 33692 40672 33744 40724
rect 33968 40715 34020 40724
rect 33968 40681 33977 40715
rect 33977 40681 34011 40715
rect 34011 40681 34020 40715
rect 33968 40672 34020 40681
rect 36176 40672 36228 40724
rect 36728 40672 36780 40724
rect 37924 40672 37976 40724
rect 34796 40647 34848 40656
rect 34796 40613 34805 40647
rect 34805 40613 34839 40647
rect 34839 40613 34848 40647
rect 34796 40604 34848 40613
rect 36544 40604 36596 40656
rect 38476 40647 38528 40656
rect 38476 40613 38485 40647
rect 38485 40613 38519 40647
rect 38519 40613 38528 40647
rect 38476 40604 38528 40613
rect 29828 40579 29880 40588
rect 29828 40545 29837 40579
rect 29837 40545 29871 40579
rect 29871 40545 29880 40579
rect 29828 40536 29880 40545
rect 30840 40536 30892 40588
rect 31668 40536 31720 40588
rect 31760 40579 31812 40588
rect 31760 40545 31769 40579
rect 31769 40545 31803 40579
rect 31803 40545 31812 40579
rect 31760 40536 31812 40545
rect 33140 40536 33192 40588
rect 36084 40536 36136 40588
rect 40500 40672 40552 40724
rect 41052 40715 41104 40724
rect 41052 40681 41061 40715
rect 41061 40681 41095 40715
rect 41095 40681 41104 40715
rect 41052 40672 41104 40681
rect 41512 40672 41564 40724
rect 42064 40715 42116 40724
rect 42064 40681 42073 40715
rect 42073 40681 42107 40715
rect 42107 40681 42116 40715
rect 42064 40672 42116 40681
rect 42248 40672 42300 40724
rect 39488 40647 39540 40656
rect 39488 40613 39497 40647
rect 39497 40613 39531 40647
rect 39531 40613 39540 40647
rect 39488 40604 39540 40613
rect 40960 40604 41012 40656
rect 42892 40604 42944 40656
rect 43168 40604 43220 40656
rect 45100 40647 45152 40656
rect 45100 40613 45109 40647
rect 45109 40613 45143 40647
rect 45143 40613 45152 40647
rect 45100 40604 45152 40613
rect 46480 40604 46532 40656
rect 47768 40647 47820 40656
rect 47768 40613 47777 40647
rect 47777 40613 47811 40647
rect 47811 40613 47820 40647
rect 47768 40604 47820 40613
rect 47952 40604 48004 40656
rect 41972 40579 42024 40588
rect 41972 40545 41981 40579
rect 41981 40545 42015 40579
rect 42015 40545 42024 40579
rect 41972 40536 42024 40545
rect 42248 40536 42300 40588
rect 47860 40579 47912 40588
rect 47860 40545 47869 40579
rect 47869 40545 47903 40579
rect 47903 40545 47912 40579
rect 47860 40536 47912 40545
rect 31116 40511 31168 40520
rect 31116 40477 31125 40511
rect 31125 40477 31159 40511
rect 31159 40477 31168 40511
rect 31116 40468 31168 40477
rect 31300 40511 31352 40520
rect 31300 40477 31309 40511
rect 31309 40477 31343 40511
rect 31343 40477 31352 40511
rect 31300 40468 31352 40477
rect 7748 40332 7800 40384
rect 15568 40332 15620 40384
rect 15752 40332 15804 40384
rect 16856 40332 16908 40384
rect 17684 40332 17736 40384
rect 17868 40375 17920 40384
rect 17868 40341 17877 40375
rect 17877 40341 17911 40375
rect 17911 40341 17920 40375
rect 17868 40332 17920 40341
rect 19340 40332 19392 40384
rect 22192 40400 22244 40452
rect 21456 40332 21508 40384
rect 21640 40332 21692 40384
rect 22008 40332 22060 40384
rect 23020 40400 23072 40452
rect 25044 40400 25096 40452
rect 27528 40400 27580 40452
rect 22744 40375 22796 40384
rect 22744 40341 22753 40375
rect 22753 40341 22787 40375
rect 22787 40341 22796 40375
rect 22744 40332 22796 40341
rect 25320 40375 25372 40384
rect 25320 40341 25329 40375
rect 25329 40341 25363 40375
rect 25363 40341 25372 40375
rect 25320 40332 25372 40341
rect 26608 40332 26660 40384
rect 29368 40375 29420 40384
rect 29368 40341 29377 40375
rect 29377 40341 29411 40375
rect 29411 40341 29420 40375
rect 29368 40332 29420 40341
rect 30564 40332 30616 40384
rect 30656 40375 30708 40384
rect 30656 40341 30665 40375
rect 30665 40341 30699 40375
rect 30699 40341 30708 40375
rect 30656 40332 30708 40341
rect 33508 40400 33560 40452
rect 34060 40511 34112 40520
rect 34060 40477 34069 40511
rect 34069 40477 34103 40511
rect 34103 40477 34112 40511
rect 34060 40468 34112 40477
rect 34152 40511 34204 40520
rect 34152 40477 34161 40511
rect 34161 40477 34195 40511
rect 34195 40477 34204 40511
rect 34152 40468 34204 40477
rect 39856 40468 39908 40520
rect 41880 40468 41932 40520
rect 44824 40511 44876 40520
rect 34888 40400 34940 40452
rect 37372 40400 37424 40452
rect 37740 40400 37792 40452
rect 41696 40400 41748 40452
rect 44824 40477 44833 40511
rect 44833 40477 44867 40511
rect 44867 40477 44876 40511
rect 44824 40468 44876 40477
rect 49700 40604 49752 40656
rect 65064 40672 65116 40724
rect 52460 40647 52512 40656
rect 52460 40613 52469 40647
rect 52469 40613 52503 40647
rect 52503 40613 52512 40647
rect 52460 40604 52512 40613
rect 53104 40604 53156 40656
rect 54024 40604 54076 40656
rect 55128 40604 55180 40656
rect 33232 40332 33284 40384
rect 34152 40332 34204 40384
rect 37096 40332 37148 40384
rect 39948 40332 40000 40384
rect 40040 40332 40092 40384
rect 42064 40332 42116 40384
rect 47216 40400 47268 40452
rect 43720 40332 43772 40384
rect 45836 40332 45888 40384
rect 49056 40511 49108 40520
rect 49056 40477 49065 40511
rect 49065 40477 49099 40511
rect 49099 40477 49108 40511
rect 49056 40468 49108 40477
rect 49148 40511 49200 40520
rect 49148 40477 49157 40511
rect 49157 40477 49191 40511
rect 49191 40477 49200 40511
rect 49148 40468 49200 40477
rect 47584 40400 47636 40452
rect 49240 40400 49292 40452
rect 48504 40332 48556 40384
rect 48596 40375 48648 40384
rect 48596 40341 48605 40375
rect 48605 40341 48639 40375
rect 48639 40341 48648 40375
rect 48596 40332 48648 40341
rect 49792 40579 49844 40588
rect 49792 40545 49801 40579
rect 49801 40545 49835 40579
rect 49835 40545 49844 40579
rect 49792 40536 49844 40545
rect 50712 40536 50764 40588
rect 52184 40579 52236 40588
rect 52184 40545 52193 40579
rect 52193 40545 52227 40579
rect 52227 40545 52236 40579
rect 52184 40536 52236 40545
rect 50436 40468 50488 40520
rect 53840 40468 53892 40520
rect 54576 40511 54628 40520
rect 54576 40477 54585 40511
rect 54585 40477 54619 40511
rect 54619 40477 54628 40511
rect 54576 40468 54628 40477
rect 55588 40468 55640 40520
rect 56048 40468 56100 40520
rect 49884 40400 49936 40452
rect 51540 40443 51592 40452
rect 51540 40409 51549 40443
rect 51549 40409 51583 40443
rect 51583 40409 51592 40443
rect 51540 40400 51592 40409
rect 50620 40332 50672 40384
rect 52644 40332 52696 40384
rect 53932 40332 53984 40384
rect 55036 40332 55088 40384
rect 1998 40230 2050 40282
rect 2062 40230 2114 40282
rect 2126 40230 2178 40282
rect 2190 40230 2242 40282
rect 2254 40230 2306 40282
rect 49998 40230 50050 40282
rect 50062 40230 50114 40282
rect 50126 40230 50178 40282
rect 50190 40230 50242 40282
rect 50254 40230 50306 40282
rect 8760 40128 8812 40180
rect 8576 40060 8628 40112
rect 9312 40035 9364 40044
rect 9312 40001 9321 40035
rect 9321 40001 9355 40035
rect 9355 40001 9364 40035
rect 9312 39992 9364 40001
rect 10508 40128 10560 40180
rect 15384 40128 15436 40180
rect 18696 40128 18748 40180
rect 10232 39992 10284 40044
rect 10968 39992 11020 40044
rect 11336 39992 11388 40044
rect 7656 39967 7708 39976
rect 7656 39933 7665 39967
rect 7665 39933 7699 39967
rect 7699 39933 7708 39967
rect 7656 39924 7708 39933
rect 12532 40060 12584 40112
rect 15476 40060 15528 40112
rect 13728 40035 13780 40044
rect 13728 40001 13737 40035
rect 13737 40001 13771 40035
rect 13771 40001 13780 40035
rect 13728 39992 13780 40001
rect 16488 39992 16540 40044
rect 18328 40060 18380 40112
rect 20720 40128 20772 40180
rect 21548 40128 21600 40180
rect 25320 40128 25372 40180
rect 27436 40128 27488 40180
rect 27528 40128 27580 40180
rect 21364 40060 21416 40112
rect 21456 40060 21508 40112
rect 12992 39924 13044 39976
rect 15476 39967 15528 39976
rect 15476 39933 15485 39967
rect 15485 39933 15519 39967
rect 15519 39933 15528 39967
rect 15476 39924 15528 39933
rect 17316 39967 17368 39976
rect 17316 39933 17325 39967
rect 17325 39933 17359 39967
rect 17359 39933 17368 39967
rect 19064 39967 19116 39976
rect 17316 39924 17368 39933
rect 19064 39933 19073 39967
rect 19073 39933 19107 39967
rect 19107 39933 19116 39967
rect 19064 39924 19116 39933
rect 20444 39924 20496 39976
rect 13912 39856 13964 39908
rect 15752 39856 15804 39908
rect 8852 39788 8904 39840
rect 9128 39831 9180 39840
rect 9128 39797 9137 39831
rect 9137 39797 9171 39831
rect 9171 39797 9180 39831
rect 9128 39788 9180 39797
rect 13084 39788 13136 39840
rect 14188 39788 14240 39840
rect 16948 39788 17000 39840
rect 17960 39831 18012 39840
rect 17960 39797 17969 39831
rect 17969 39797 18003 39831
rect 18003 39797 18012 39831
rect 17960 39788 18012 39797
rect 18144 39788 18196 39840
rect 21272 39967 21324 39976
rect 21272 39933 21281 39967
rect 21281 39933 21315 39967
rect 21315 39933 21324 39967
rect 21272 39924 21324 39933
rect 21824 39992 21876 40044
rect 22284 40035 22336 40044
rect 22284 40001 22293 40035
rect 22293 40001 22327 40035
rect 22327 40001 22336 40035
rect 22284 39992 22336 40001
rect 22928 40060 22980 40112
rect 29828 40128 29880 40180
rect 30656 40128 30708 40180
rect 31484 40171 31536 40180
rect 31484 40137 31493 40171
rect 31493 40137 31527 40171
rect 31527 40137 31536 40171
rect 31484 40128 31536 40137
rect 33048 40171 33100 40180
rect 33048 40137 33069 40171
rect 33069 40137 33100 40171
rect 33048 40128 33100 40137
rect 34060 40128 34112 40180
rect 37464 40128 37516 40180
rect 38108 40128 38160 40180
rect 39672 40128 39724 40180
rect 41420 40128 41472 40180
rect 22652 40035 22704 40044
rect 22652 40001 22661 40035
rect 22661 40001 22695 40035
rect 22695 40001 22704 40035
rect 22652 39992 22704 40001
rect 23296 40035 23348 40044
rect 23296 40001 23305 40035
rect 23305 40001 23339 40035
rect 23339 40001 23348 40035
rect 23296 39992 23348 40001
rect 26516 39992 26568 40044
rect 27160 39992 27212 40044
rect 33508 40060 33560 40112
rect 34520 40060 34572 40112
rect 31852 39992 31904 40044
rect 23480 39924 23532 39976
rect 24032 39924 24084 39976
rect 26240 39924 26292 39976
rect 29552 39924 29604 39976
rect 32588 39992 32640 40044
rect 34980 40060 35032 40112
rect 39396 40060 39448 40112
rect 37280 39992 37332 40044
rect 37372 40035 37424 40044
rect 37372 40001 37381 40035
rect 37381 40001 37415 40035
rect 37415 40001 37424 40035
rect 37372 39992 37424 40001
rect 38660 39992 38712 40044
rect 41604 40060 41656 40112
rect 43352 40128 43404 40180
rect 45744 40128 45796 40180
rect 21732 39856 21784 39908
rect 24860 39856 24912 39908
rect 24952 39856 25004 39908
rect 21272 39788 21324 39840
rect 23848 39831 23900 39840
rect 23848 39797 23857 39831
rect 23857 39797 23891 39831
rect 23891 39797 23900 39831
rect 23848 39788 23900 39797
rect 32588 39856 32640 39908
rect 32956 39856 33008 39908
rect 33784 39856 33836 39908
rect 34888 39924 34940 39976
rect 39764 39967 39816 39976
rect 39764 39933 39773 39967
rect 39773 39933 39807 39967
rect 39807 39933 39816 39967
rect 39764 39924 39816 39933
rect 41052 39924 41104 39976
rect 35624 39856 35676 39908
rect 36084 39856 36136 39908
rect 38108 39856 38160 39908
rect 40040 39899 40092 39908
rect 40040 39865 40049 39899
rect 40049 39865 40083 39899
rect 40083 39865 40092 39899
rect 40040 39856 40092 39865
rect 43812 40060 43864 40112
rect 43076 40035 43128 40044
rect 43076 40001 43085 40035
rect 43085 40001 43119 40035
rect 43119 40001 43128 40035
rect 43076 39992 43128 40001
rect 43536 39992 43588 40044
rect 43996 40060 44048 40112
rect 44824 40035 44876 40044
rect 44824 40001 44833 40035
rect 44833 40001 44867 40035
rect 44867 40001 44876 40035
rect 44824 39992 44876 40001
rect 46112 39992 46164 40044
rect 48596 40128 48648 40180
rect 49608 40128 49660 40180
rect 51356 40128 51408 40180
rect 49884 40060 49936 40112
rect 50436 40060 50488 40112
rect 49700 40035 49752 40044
rect 49700 40001 49709 40035
rect 49709 40001 49743 40035
rect 49743 40001 49752 40035
rect 49700 39992 49752 40001
rect 42156 39924 42208 39976
rect 26332 39831 26384 39840
rect 26332 39797 26341 39831
rect 26341 39797 26375 39831
rect 26375 39797 26384 39831
rect 26332 39788 26384 39797
rect 27068 39788 27120 39840
rect 27436 39788 27488 39840
rect 28356 39788 28408 39840
rect 31024 39788 31076 39840
rect 41052 39788 41104 39840
rect 41512 39831 41564 39840
rect 41512 39797 41521 39831
rect 41521 39797 41555 39831
rect 41555 39797 41564 39831
rect 41512 39788 41564 39797
rect 41604 39831 41656 39840
rect 41604 39797 41613 39831
rect 41613 39797 41647 39831
rect 41647 39797 41656 39831
rect 41604 39788 41656 39797
rect 41972 39788 42024 39840
rect 43536 39788 43588 39840
rect 43720 39831 43772 39840
rect 43720 39797 43729 39831
rect 43729 39797 43763 39831
rect 43763 39797 43772 39831
rect 43720 39788 43772 39797
rect 46480 39856 46532 39908
rect 46664 39831 46716 39840
rect 46664 39797 46673 39831
rect 46673 39797 46707 39831
rect 46707 39797 46716 39831
rect 46664 39788 46716 39797
rect 48964 39856 49016 39908
rect 49884 39831 49936 39840
rect 49884 39797 49893 39831
rect 49893 39797 49927 39831
rect 49927 39797 49936 39831
rect 49884 39788 49936 39797
rect 49976 39831 50028 39840
rect 49976 39797 49985 39831
rect 49985 39797 50019 39831
rect 50019 39797 50028 39831
rect 49976 39788 50028 39797
rect 50252 39788 50304 39840
rect 50712 39899 50764 39908
rect 50712 39865 50721 39899
rect 50721 39865 50755 39899
rect 50755 39865 50764 39899
rect 51540 40060 51592 40112
rect 53472 39992 53524 40044
rect 54576 40128 54628 40180
rect 55588 40171 55640 40180
rect 55588 40137 55597 40171
rect 55597 40137 55631 40171
rect 55631 40137 55640 40171
rect 55588 40128 55640 40137
rect 55036 40060 55088 40112
rect 60740 40060 60792 40112
rect 64972 40060 65024 40112
rect 54668 39992 54720 40044
rect 56232 40035 56284 40044
rect 56232 40001 56241 40035
rect 56241 40001 56275 40035
rect 56275 40001 56284 40035
rect 56232 39992 56284 40001
rect 56508 39924 56560 39976
rect 50712 39856 50764 39865
rect 52092 39899 52144 39908
rect 52092 39865 52101 39899
rect 52101 39865 52135 39899
rect 52135 39865 52144 39899
rect 52092 39856 52144 39865
rect 53104 39856 53156 39908
rect 56048 39899 56100 39908
rect 52828 39788 52880 39840
rect 54484 39788 54536 39840
rect 56048 39865 56057 39899
rect 56057 39865 56091 39899
rect 56091 39865 56100 39899
rect 56048 39856 56100 39865
rect 55312 39788 55364 39840
rect 2918 39686 2970 39738
rect 2982 39686 3034 39738
rect 3046 39686 3098 39738
rect 3110 39686 3162 39738
rect 3174 39686 3226 39738
rect 50918 39686 50970 39738
rect 50982 39686 51034 39738
rect 51046 39686 51098 39738
rect 51110 39686 51162 39738
rect 51174 39686 51226 39738
rect 8576 39516 8628 39568
rect 8852 39559 8904 39568
rect 8852 39525 8861 39559
rect 8861 39525 8895 39559
rect 8895 39525 8904 39559
rect 8852 39516 8904 39525
rect 12808 39584 12860 39636
rect 9496 39516 9548 39568
rect 11428 39559 11480 39568
rect 11428 39525 11437 39559
rect 11437 39525 11471 39559
rect 11471 39525 11480 39559
rect 11428 39516 11480 39525
rect 12440 39516 12492 39568
rect 13544 39516 13596 39568
rect 7656 39380 7708 39432
rect 11704 39448 11756 39500
rect 15476 39516 15528 39568
rect 15568 39559 15620 39568
rect 15568 39525 15577 39559
rect 15577 39525 15611 39559
rect 15611 39525 15620 39559
rect 15568 39516 15620 39525
rect 13912 39448 13964 39500
rect 14464 39448 14516 39500
rect 17316 39584 17368 39636
rect 18420 39627 18472 39636
rect 18420 39593 18429 39627
rect 18429 39593 18463 39627
rect 18463 39593 18472 39627
rect 18420 39584 18472 39593
rect 19064 39584 19116 39636
rect 21272 39627 21324 39636
rect 21272 39593 21281 39627
rect 21281 39593 21315 39627
rect 21315 39593 21324 39627
rect 21272 39584 21324 39593
rect 21364 39584 21416 39636
rect 22744 39584 22796 39636
rect 24032 39627 24084 39636
rect 24032 39593 24041 39627
rect 24041 39593 24075 39627
rect 24075 39593 24084 39627
rect 24032 39584 24084 39593
rect 25136 39627 25188 39636
rect 25136 39593 25145 39627
rect 25145 39593 25179 39627
rect 25179 39593 25188 39627
rect 25136 39584 25188 39593
rect 26332 39584 26384 39636
rect 16948 39559 17000 39568
rect 16948 39525 16957 39559
rect 16957 39525 16991 39559
rect 16991 39525 17000 39559
rect 16948 39516 17000 39525
rect 18512 39516 18564 39568
rect 24676 39516 24728 39568
rect 24860 39516 24912 39568
rect 28356 39584 28408 39636
rect 28724 39584 28776 39636
rect 29368 39584 29420 39636
rect 31484 39584 31536 39636
rect 27620 39516 27672 39568
rect 30380 39516 30432 39568
rect 33232 39584 33284 39636
rect 33600 39584 33652 39636
rect 33692 39584 33744 39636
rect 34612 39584 34664 39636
rect 35256 39584 35308 39636
rect 35992 39584 36044 39636
rect 18052 39448 18104 39500
rect 21548 39448 21600 39500
rect 21732 39491 21784 39500
rect 21732 39457 21741 39491
rect 21741 39457 21775 39491
rect 21775 39457 21784 39491
rect 21732 39448 21784 39457
rect 9588 39312 9640 39364
rect 13084 39380 13136 39432
rect 10416 39312 10468 39364
rect 14372 39423 14424 39432
rect 14372 39389 14381 39423
rect 14381 39389 14415 39423
rect 14415 39389 14424 39423
rect 14372 39380 14424 39389
rect 15292 39423 15344 39432
rect 15292 39389 15301 39423
rect 15301 39389 15335 39423
rect 15335 39389 15344 39423
rect 15292 39380 15344 39389
rect 17408 39380 17460 39432
rect 20812 39380 20864 39432
rect 21824 39423 21876 39432
rect 21824 39389 21833 39423
rect 21833 39389 21867 39423
rect 21867 39389 21876 39423
rect 21824 39380 21876 39389
rect 15936 39355 15988 39364
rect 15936 39321 15945 39355
rect 15945 39321 15979 39355
rect 15979 39321 15988 39355
rect 15936 39312 15988 39321
rect 8852 39244 8904 39296
rect 12992 39244 13044 39296
rect 20536 39244 20588 39296
rect 22652 39423 22704 39432
rect 22652 39389 22661 39423
rect 22661 39389 22695 39423
rect 22695 39389 22704 39423
rect 22652 39380 22704 39389
rect 22468 39312 22520 39364
rect 24308 39380 24360 39432
rect 25596 39423 25648 39432
rect 25596 39389 25605 39423
rect 25605 39389 25639 39423
rect 25639 39389 25648 39423
rect 25596 39380 25648 39389
rect 28724 39448 28776 39500
rect 26424 39380 26476 39432
rect 26056 39312 26108 39364
rect 27620 39312 27672 39364
rect 28816 39380 28868 39432
rect 34520 39516 34572 39568
rect 29000 39423 29052 39432
rect 29000 39389 29009 39423
rect 29009 39389 29043 39423
rect 29043 39389 29052 39423
rect 29000 39380 29052 39389
rect 27896 39312 27948 39364
rect 31576 39491 31628 39500
rect 31576 39457 31585 39491
rect 31585 39457 31619 39491
rect 31619 39457 31628 39491
rect 31576 39448 31628 39457
rect 32956 39448 33008 39500
rect 33416 39448 33468 39500
rect 36636 39516 36688 39568
rect 37004 39559 37056 39568
rect 37004 39525 37013 39559
rect 37013 39525 37047 39559
rect 37047 39525 37056 39559
rect 37004 39516 37056 39525
rect 38568 39627 38620 39636
rect 38568 39593 38577 39627
rect 38577 39593 38611 39627
rect 38611 39593 38620 39627
rect 38568 39584 38620 39593
rect 38936 39627 38988 39636
rect 38936 39593 38945 39627
rect 38945 39593 38979 39627
rect 38979 39593 38988 39627
rect 38936 39584 38988 39593
rect 36544 39448 36596 39500
rect 36728 39491 36780 39500
rect 36728 39457 36737 39491
rect 36737 39457 36771 39491
rect 36771 39457 36780 39491
rect 36728 39448 36780 39457
rect 38108 39448 38160 39500
rect 40960 39516 41012 39568
rect 42984 39584 43036 39636
rect 44088 39584 44140 39636
rect 46112 39627 46164 39636
rect 46112 39593 46121 39627
rect 46121 39593 46155 39627
rect 46155 39593 46164 39627
rect 46112 39584 46164 39593
rect 46664 39584 46716 39636
rect 48412 39584 48464 39636
rect 49884 39584 49936 39636
rect 49976 39584 50028 39636
rect 41512 39516 41564 39568
rect 43444 39516 43496 39568
rect 45744 39516 45796 39568
rect 42432 39491 42484 39500
rect 42432 39457 42441 39491
rect 42441 39457 42475 39491
rect 42475 39457 42484 39491
rect 42432 39448 42484 39457
rect 42708 39448 42760 39500
rect 30104 39380 30156 39432
rect 30840 39380 30892 39432
rect 24124 39244 24176 39296
rect 25964 39244 26016 39296
rect 26516 39244 26568 39296
rect 27252 39244 27304 39296
rect 29000 39244 29052 39296
rect 29092 39244 29144 39296
rect 32220 39380 32272 39432
rect 32588 39380 32640 39432
rect 37372 39380 37424 39432
rect 37464 39380 37516 39432
rect 38568 39380 38620 39432
rect 39120 39423 39172 39432
rect 39120 39389 39129 39423
rect 39129 39389 39163 39423
rect 39163 39389 39172 39423
rect 39120 39380 39172 39389
rect 33232 39312 33284 39364
rect 32404 39244 32456 39296
rect 33508 39244 33560 39296
rect 35624 39312 35676 39364
rect 36728 39312 36780 39364
rect 41420 39380 41472 39432
rect 41788 39380 41840 39432
rect 41880 39380 41932 39432
rect 42616 39423 42668 39432
rect 42616 39389 42625 39423
rect 42625 39389 42659 39423
rect 42659 39389 42668 39423
rect 42616 39380 42668 39389
rect 37464 39244 37516 39296
rect 37556 39244 37608 39296
rect 38752 39244 38804 39296
rect 40408 39312 40460 39364
rect 40132 39244 40184 39296
rect 41052 39244 41104 39296
rect 41972 39312 42024 39364
rect 42156 39312 42208 39364
rect 43444 39423 43496 39432
rect 43444 39389 43453 39423
rect 43453 39389 43487 39423
rect 43487 39389 43496 39423
rect 43444 39380 43496 39389
rect 45284 39448 45336 39500
rect 45100 39423 45152 39432
rect 45100 39389 45109 39423
rect 45109 39389 45143 39423
rect 45143 39389 45152 39423
rect 45836 39448 45888 39500
rect 46020 39516 46072 39568
rect 46296 39448 46348 39500
rect 48320 39516 48372 39568
rect 48872 39516 48924 39568
rect 50252 39559 50304 39568
rect 50252 39525 50261 39559
rect 50261 39525 50295 39559
rect 50295 39525 50304 39559
rect 50252 39516 50304 39525
rect 50620 39559 50672 39568
rect 50620 39525 50629 39559
rect 50629 39525 50663 39559
rect 50663 39525 50672 39559
rect 50620 39516 50672 39525
rect 48780 39448 48832 39500
rect 52368 39627 52420 39636
rect 52368 39593 52377 39627
rect 52377 39593 52411 39627
rect 52411 39593 52420 39627
rect 52368 39584 52420 39593
rect 52736 39584 52788 39636
rect 63500 39584 63552 39636
rect 51356 39559 51408 39568
rect 51356 39525 51365 39559
rect 51365 39525 51399 39559
rect 51399 39525 51408 39559
rect 51356 39516 51408 39525
rect 52184 39516 52236 39568
rect 52828 39559 52880 39568
rect 52828 39525 52837 39559
rect 52837 39525 52871 39559
rect 52871 39525 52880 39559
rect 52828 39516 52880 39525
rect 54760 39516 54812 39568
rect 52092 39448 52144 39500
rect 52644 39448 52696 39500
rect 45100 39380 45152 39389
rect 45560 39423 45612 39432
rect 45560 39389 45569 39423
rect 45569 39389 45603 39423
rect 45603 39389 45612 39423
rect 45560 39380 45612 39389
rect 45928 39312 45980 39364
rect 46756 39423 46808 39432
rect 46756 39389 46765 39423
rect 46765 39389 46799 39423
rect 46799 39389 46808 39423
rect 46756 39380 46808 39389
rect 41788 39244 41840 39296
rect 42340 39244 42392 39296
rect 48412 39380 48464 39432
rect 48136 39312 48188 39364
rect 50712 39380 50764 39432
rect 54668 39448 54720 39500
rect 59268 39516 59320 39568
rect 53564 39380 53616 39432
rect 55956 39423 56008 39432
rect 55956 39389 55965 39423
rect 55965 39389 55999 39423
rect 55999 39389 56008 39423
rect 55956 39380 56008 39389
rect 56324 39380 56376 39432
rect 56784 39380 56836 39432
rect 50804 39312 50856 39364
rect 56692 39312 56744 39364
rect 59912 39312 59964 39364
rect 47400 39244 47452 39296
rect 53196 39287 53248 39296
rect 53196 39253 53205 39287
rect 53205 39253 53239 39287
rect 53239 39253 53248 39287
rect 53196 39244 53248 39253
rect 55312 39244 55364 39296
rect 56232 39244 56284 39296
rect 59176 39244 59228 39296
rect 60280 39287 60332 39296
rect 60280 39253 60289 39287
rect 60289 39253 60323 39287
rect 60323 39253 60332 39287
rect 60280 39244 60332 39253
rect 60372 39287 60424 39296
rect 60372 39253 60381 39287
rect 60381 39253 60415 39287
rect 60415 39253 60424 39287
rect 60372 39244 60424 39253
rect 1998 39142 2050 39194
rect 2062 39142 2114 39194
rect 2126 39142 2178 39194
rect 2190 39142 2242 39194
rect 2254 39142 2306 39194
rect 49998 39142 50050 39194
rect 50062 39142 50114 39194
rect 50126 39142 50178 39194
rect 50190 39142 50242 39194
rect 50254 39142 50306 39194
rect 8576 39040 8628 39092
rect 8760 38904 8812 38956
rect 8668 38768 8720 38820
rect 8852 38768 8904 38820
rect 11428 39040 11480 39092
rect 11520 38904 11572 38956
rect 7564 38743 7616 38752
rect 7564 38709 7573 38743
rect 7573 38709 7607 38743
rect 7607 38709 7616 38743
rect 7564 38700 7616 38709
rect 10876 38811 10928 38820
rect 10876 38777 10885 38811
rect 10885 38777 10919 38811
rect 10919 38777 10928 38811
rect 10876 38768 10928 38777
rect 10968 38768 11020 38820
rect 12808 38947 12860 38956
rect 12808 38913 12817 38947
rect 12817 38913 12851 38947
rect 12851 38913 12860 38947
rect 12808 38904 12860 38913
rect 20168 39040 20220 39092
rect 23940 39040 23992 39092
rect 24308 39040 24360 39092
rect 26056 39040 26108 39092
rect 15200 38972 15252 39024
rect 16396 38972 16448 39024
rect 21732 38972 21784 39024
rect 25596 39015 25648 39024
rect 25596 38981 25605 39015
rect 25605 38981 25639 39015
rect 25639 38981 25648 39015
rect 25596 38972 25648 38981
rect 26700 38972 26752 39024
rect 13820 38904 13872 38956
rect 14832 38904 14884 38956
rect 16764 38947 16816 38956
rect 16764 38913 16773 38947
rect 16773 38913 16807 38947
rect 16807 38913 16816 38947
rect 16764 38904 16816 38913
rect 19064 38904 19116 38956
rect 21916 38947 21968 38956
rect 21916 38913 21925 38947
rect 21925 38913 21959 38947
rect 21959 38913 21968 38947
rect 21916 38904 21968 38913
rect 22192 38904 22244 38956
rect 23388 38904 23440 38956
rect 24124 38947 24176 38956
rect 24124 38913 24133 38947
rect 24133 38913 24167 38947
rect 24167 38913 24176 38947
rect 24124 38904 24176 38913
rect 24216 38904 24268 38956
rect 24492 38904 24544 38956
rect 27988 39040 28040 39092
rect 42340 39040 42392 39092
rect 42432 39040 42484 39092
rect 45284 39083 45336 39092
rect 45284 39049 45293 39083
rect 45293 39049 45327 39083
rect 45327 39049 45336 39083
rect 45284 39040 45336 39049
rect 46020 39040 46072 39092
rect 49056 39040 49108 39092
rect 30104 38904 30156 38956
rect 30288 38904 30340 38956
rect 12992 38879 13044 38888
rect 12992 38845 13001 38879
rect 13001 38845 13035 38879
rect 13035 38845 13044 38879
rect 12992 38836 13044 38845
rect 15292 38836 15344 38888
rect 21732 38879 21784 38888
rect 21732 38845 21741 38879
rect 21741 38845 21775 38879
rect 21775 38845 21784 38879
rect 21732 38836 21784 38845
rect 26516 38836 26568 38888
rect 26700 38836 26752 38888
rect 30472 38904 30524 38956
rect 31116 38972 31168 39024
rect 33600 38972 33652 39024
rect 32220 38947 32272 38956
rect 32220 38913 32229 38947
rect 32229 38913 32263 38947
rect 32263 38913 32272 38947
rect 32220 38904 32272 38913
rect 31668 38836 31720 38888
rect 32404 38879 32456 38888
rect 32404 38845 32413 38879
rect 32413 38845 32447 38879
rect 32447 38845 32456 38879
rect 32404 38836 32456 38845
rect 13452 38768 13504 38820
rect 12348 38743 12400 38752
rect 12348 38709 12357 38743
rect 12357 38709 12391 38743
rect 12391 38709 12400 38743
rect 12348 38700 12400 38709
rect 14096 38768 14148 38820
rect 19524 38768 19576 38820
rect 19616 38811 19668 38820
rect 19616 38777 19625 38811
rect 19625 38777 19659 38811
rect 19659 38777 19668 38811
rect 19616 38768 19668 38777
rect 15384 38700 15436 38752
rect 18052 38700 18104 38752
rect 19248 38700 19300 38752
rect 22192 38811 22244 38820
rect 22192 38777 22201 38811
rect 22201 38777 22235 38811
rect 22235 38777 22244 38811
rect 22192 38768 22244 38777
rect 21364 38700 21416 38752
rect 22008 38700 22060 38752
rect 28908 38768 28960 38820
rect 29000 38768 29052 38820
rect 24952 38700 25004 38752
rect 25688 38743 25740 38752
rect 25688 38709 25697 38743
rect 25697 38709 25731 38743
rect 25731 38709 25740 38743
rect 25688 38700 25740 38709
rect 26148 38743 26200 38752
rect 26148 38709 26157 38743
rect 26157 38709 26191 38743
rect 26191 38709 26200 38743
rect 26148 38700 26200 38709
rect 26792 38700 26844 38752
rect 27712 38700 27764 38752
rect 27804 38700 27856 38752
rect 28264 38743 28316 38752
rect 28264 38709 28273 38743
rect 28273 38709 28307 38743
rect 28307 38709 28316 38743
rect 28264 38700 28316 38709
rect 29092 38700 29144 38752
rect 29184 38700 29236 38752
rect 29920 38743 29972 38752
rect 29920 38709 29929 38743
rect 29929 38709 29963 38743
rect 29963 38709 29972 38743
rect 29920 38700 29972 38709
rect 30656 38768 30708 38820
rect 31944 38811 31996 38820
rect 31944 38777 31953 38811
rect 31953 38777 31987 38811
rect 31987 38777 31996 38811
rect 33968 38879 34020 38888
rect 33968 38845 33977 38879
rect 33977 38845 34011 38879
rect 34011 38845 34020 38879
rect 33968 38836 34020 38845
rect 31944 38768 31996 38777
rect 33232 38768 33284 38820
rect 33508 38768 33560 38820
rect 33784 38768 33836 38820
rect 35624 38947 35676 38956
rect 35624 38913 35633 38947
rect 35633 38913 35667 38947
rect 35667 38913 35676 38947
rect 35624 38904 35676 38913
rect 37556 38972 37608 39024
rect 37648 39015 37700 39024
rect 37648 38981 37657 39015
rect 37657 38981 37691 39015
rect 37691 38981 37700 39015
rect 37648 38972 37700 38981
rect 37740 38972 37792 39024
rect 37372 38904 37424 38956
rect 34704 38700 34756 38752
rect 34888 38743 34940 38752
rect 34888 38709 34897 38743
rect 34897 38709 34931 38743
rect 34931 38709 34940 38743
rect 34888 38700 34940 38709
rect 37280 38836 37332 38888
rect 38292 38836 38344 38888
rect 39212 38972 39264 39024
rect 39396 38972 39448 39024
rect 40132 38972 40184 39024
rect 40408 38972 40460 39024
rect 39488 38904 39540 38956
rect 40500 38904 40552 38956
rect 40684 38947 40736 38956
rect 40684 38913 40693 38947
rect 40693 38913 40727 38947
rect 40727 38913 40736 38947
rect 40684 38904 40736 38913
rect 40960 38904 41012 38956
rect 41328 38904 41380 38956
rect 39580 38836 39632 38888
rect 39764 38836 39816 38888
rect 42524 38904 42576 38956
rect 43260 38947 43312 38956
rect 43260 38913 43269 38947
rect 43269 38913 43303 38947
rect 43303 38913 43312 38947
rect 43260 38904 43312 38913
rect 44364 38904 44416 38956
rect 47124 38904 47176 38956
rect 48688 38904 48740 38956
rect 49240 38947 49292 38956
rect 49240 38913 49249 38947
rect 49249 38913 49283 38947
rect 49283 38913 49292 38947
rect 49240 38904 49292 38913
rect 56048 38904 56100 38956
rect 56324 38904 56376 38956
rect 57428 38904 57480 38956
rect 60464 39040 60516 39092
rect 59544 38972 59596 39024
rect 59176 38904 59228 38956
rect 59636 38904 59688 38956
rect 43720 38836 43772 38888
rect 46480 38836 46532 38888
rect 47860 38879 47912 38888
rect 47860 38845 47869 38879
rect 47869 38845 47903 38879
rect 47903 38845 47912 38879
rect 47860 38836 47912 38845
rect 48136 38836 48188 38888
rect 48412 38836 48464 38888
rect 51448 38879 51500 38888
rect 51448 38845 51457 38879
rect 51457 38845 51491 38879
rect 51491 38845 51500 38879
rect 51448 38836 51500 38845
rect 57796 38836 57848 38888
rect 60280 38836 60332 38888
rect 35900 38811 35952 38820
rect 35900 38777 35909 38811
rect 35909 38777 35943 38811
rect 35943 38777 35952 38811
rect 35900 38768 35952 38777
rect 37188 38768 37240 38820
rect 37464 38811 37516 38820
rect 37464 38777 37473 38811
rect 37473 38777 37507 38811
rect 37507 38777 37516 38811
rect 37464 38768 37516 38777
rect 36820 38700 36872 38752
rect 37372 38743 37424 38752
rect 37372 38709 37381 38743
rect 37381 38709 37415 38743
rect 37415 38709 37424 38743
rect 37372 38700 37424 38709
rect 39120 38743 39172 38752
rect 39120 38709 39129 38743
rect 39129 38709 39163 38743
rect 39163 38709 39172 38743
rect 39120 38700 39172 38709
rect 41788 38811 41840 38820
rect 41788 38777 41797 38811
rect 41797 38777 41831 38811
rect 41831 38777 41840 38811
rect 41788 38768 41840 38777
rect 40132 38743 40184 38752
rect 40132 38709 40141 38743
rect 40141 38709 40175 38743
rect 40175 38709 40184 38743
rect 40132 38700 40184 38709
rect 40500 38743 40552 38752
rect 40500 38709 40509 38743
rect 40509 38709 40543 38743
rect 40543 38709 40552 38743
rect 40500 38700 40552 38709
rect 41052 38700 41104 38752
rect 45652 38768 45704 38820
rect 47584 38811 47636 38820
rect 47584 38777 47593 38811
rect 47593 38777 47627 38811
rect 47627 38777 47636 38811
rect 47584 38768 47636 38777
rect 53012 38768 53064 38820
rect 53656 38811 53708 38820
rect 53656 38777 53665 38811
rect 53665 38777 53699 38811
rect 53699 38777 53708 38811
rect 53656 38768 53708 38777
rect 55312 38811 55364 38820
rect 55312 38777 55321 38811
rect 55321 38777 55355 38811
rect 55355 38777 55364 38811
rect 55312 38768 55364 38777
rect 44088 38700 44140 38752
rect 44916 38743 44968 38752
rect 44916 38709 44925 38743
rect 44925 38709 44959 38743
rect 44959 38709 44968 38743
rect 44916 38700 44968 38709
rect 46940 38700 46992 38752
rect 47860 38700 47912 38752
rect 49884 38743 49936 38752
rect 49884 38709 49893 38743
rect 49893 38709 49927 38743
rect 49927 38709 49936 38743
rect 49884 38700 49936 38709
rect 50344 38743 50396 38752
rect 50344 38709 50353 38743
rect 50353 38709 50387 38743
rect 50387 38709 50396 38743
rect 50344 38700 50396 38709
rect 53564 38700 53616 38752
rect 55220 38700 55272 38752
rect 55772 38768 55824 38820
rect 56784 38743 56836 38752
rect 56784 38709 56793 38743
rect 56793 38709 56827 38743
rect 56827 38709 56836 38743
rect 56784 38700 56836 38709
rect 58164 38700 58216 38752
rect 59176 38700 59228 38752
rect 2918 38598 2970 38650
rect 2982 38598 3034 38650
rect 3046 38598 3098 38650
rect 3110 38598 3162 38650
rect 3174 38598 3226 38650
rect 50918 38598 50970 38650
rect 50982 38598 51034 38650
rect 51046 38598 51098 38650
rect 51110 38598 51162 38650
rect 51174 38598 51226 38650
rect 8392 38496 8444 38548
rect 8668 38496 8720 38548
rect 8852 38539 8904 38548
rect 8852 38505 8861 38539
rect 8861 38505 8895 38539
rect 8895 38505 8904 38539
rect 8852 38496 8904 38505
rect 9128 38496 9180 38548
rect 9496 38496 9548 38548
rect 10876 38496 10928 38548
rect 11244 38496 11296 38548
rect 9956 38360 10008 38412
rect 7472 38292 7524 38344
rect 9680 38335 9732 38344
rect 9680 38301 9689 38335
rect 9689 38301 9723 38335
rect 9723 38301 9732 38335
rect 9680 38292 9732 38301
rect 11244 38360 11296 38412
rect 12348 38360 12400 38412
rect 13636 38496 13688 38548
rect 14464 38539 14516 38548
rect 14464 38505 14473 38539
rect 14473 38505 14507 38539
rect 14507 38505 14516 38539
rect 14464 38496 14516 38505
rect 16488 38496 16540 38548
rect 19340 38496 19392 38548
rect 20536 38539 20588 38548
rect 20536 38505 20545 38539
rect 20545 38505 20579 38539
rect 20579 38505 20588 38539
rect 20536 38496 20588 38505
rect 21640 38539 21692 38548
rect 21640 38505 21649 38539
rect 21649 38505 21683 38539
rect 21683 38505 21692 38539
rect 21640 38496 21692 38505
rect 15200 38428 15252 38480
rect 15476 38428 15528 38480
rect 19248 38428 19300 38480
rect 22100 38496 22152 38548
rect 22192 38496 22244 38548
rect 23848 38496 23900 38548
rect 24584 38496 24636 38548
rect 21916 38428 21968 38480
rect 9312 38224 9364 38276
rect 11336 38292 11388 38344
rect 12808 38292 12860 38344
rect 13728 38292 13780 38344
rect 15292 38360 15344 38412
rect 10968 38156 11020 38208
rect 12624 38224 12676 38276
rect 14556 38224 14608 38276
rect 16488 38403 16540 38412
rect 16488 38369 16497 38403
rect 16497 38369 16531 38403
rect 16531 38369 16540 38403
rect 16488 38360 16540 38369
rect 17592 38403 17644 38412
rect 17592 38369 17601 38403
rect 17601 38369 17635 38403
rect 17635 38369 17644 38403
rect 17592 38360 17644 38369
rect 17684 38360 17736 38412
rect 16396 38292 16448 38344
rect 18788 38292 18840 38344
rect 14372 38156 14424 38208
rect 15200 38199 15252 38208
rect 15200 38165 15209 38199
rect 15209 38165 15243 38199
rect 15243 38165 15252 38199
rect 15200 38156 15252 38165
rect 17868 38224 17920 38276
rect 19248 38156 19300 38208
rect 19340 38156 19392 38208
rect 20720 38224 20772 38276
rect 21456 38224 21508 38276
rect 21732 38335 21784 38344
rect 21732 38301 21741 38335
rect 21741 38301 21775 38335
rect 21775 38301 21784 38335
rect 21732 38292 21784 38301
rect 20904 38156 20956 38208
rect 22468 38403 22520 38412
rect 22468 38369 22477 38403
rect 22477 38369 22511 38403
rect 22511 38369 22520 38403
rect 22468 38360 22520 38369
rect 25044 38428 25096 38480
rect 26240 38496 26292 38548
rect 26976 38428 27028 38480
rect 27620 38428 27672 38480
rect 28448 38360 28500 38412
rect 29552 38496 29604 38548
rect 29920 38496 29972 38548
rect 33140 38496 33192 38548
rect 29184 38471 29236 38480
rect 29184 38437 29193 38471
rect 29193 38437 29227 38471
rect 29227 38437 29236 38471
rect 29184 38428 29236 38437
rect 31208 38428 31260 38480
rect 31392 38428 31444 38480
rect 33876 38428 33928 38480
rect 34888 38496 34940 38548
rect 35900 38496 35952 38548
rect 36820 38496 36872 38548
rect 38292 38496 38344 38548
rect 23572 38335 23624 38344
rect 23572 38301 23581 38335
rect 23581 38301 23615 38335
rect 23615 38301 23624 38335
rect 23572 38292 23624 38301
rect 24032 38292 24084 38344
rect 25688 38292 25740 38344
rect 27068 38335 27120 38344
rect 27068 38301 27077 38335
rect 27077 38301 27111 38335
rect 27111 38301 27120 38335
rect 27068 38292 27120 38301
rect 30748 38292 30800 38344
rect 32956 38360 33008 38412
rect 33232 38360 33284 38412
rect 34888 38403 34940 38412
rect 34888 38369 34897 38403
rect 34897 38369 34931 38403
rect 34931 38369 34940 38403
rect 34888 38360 34940 38369
rect 36268 38471 36320 38480
rect 36268 38437 36277 38471
rect 36277 38437 36311 38471
rect 36311 38437 36320 38471
rect 36268 38428 36320 38437
rect 37372 38360 37424 38412
rect 28356 38224 28408 38276
rect 25872 38199 25924 38208
rect 25872 38165 25881 38199
rect 25881 38165 25915 38199
rect 25915 38165 25924 38199
rect 25872 38156 25924 38165
rect 27528 38156 27580 38208
rect 28816 38199 28868 38208
rect 28816 38165 28825 38199
rect 28825 38165 28859 38199
rect 28859 38165 28868 38199
rect 28816 38156 28868 38165
rect 32956 38156 33008 38208
rect 33232 38156 33284 38208
rect 34888 38224 34940 38276
rect 35164 38292 35216 38344
rect 35440 38292 35492 38344
rect 35716 38292 35768 38344
rect 39212 38428 39264 38480
rect 39672 38428 39724 38480
rect 40040 38496 40092 38548
rect 41236 38496 41288 38548
rect 42524 38496 42576 38548
rect 40224 38428 40276 38480
rect 41144 38428 41196 38480
rect 43444 38471 43496 38480
rect 43444 38437 43453 38471
rect 43453 38437 43487 38471
rect 43487 38437 43496 38471
rect 43444 38428 43496 38437
rect 41236 38360 41288 38412
rect 41328 38360 41380 38412
rect 44824 38496 44876 38548
rect 45652 38539 45704 38548
rect 45652 38505 45661 38539
rect 45661 38505 45695 38539
rect 45695 38505 45704 38539
rect 45652 38496 45704 38505
rect 47400 38539 47452 38548
rect 47400 38505 47409 38539
rect 47409 38505 47443 38539
rect 47443 38505 47452 38539
rect 47400 38496 47452 38505
rect 47584 38496 47636 38548
rect 48688 38496 48740 38548
rect 48780 38539 48832 38548
rect 48780 38505 48789 38539
rect 48789 38505 48823 38539
rect 48823 38505 48832 38539
rect 48780 38496 48832 38505
rect 51448 38496 51500 38548
rect 53196 38496 53248 38548
rect 53656 38539 53708 38548
rect 53656 38505 53665 38539
rect 53665 38505 53699 38539
rect 53699 38505 53708 38539
rect 53656 38496 53708 38505
rect 44088 38471 44140 38480
rect 44088 38437 44097 38471
rect 44097 38437 44131 38471
rect 44131 38437 44140 38471
rect 44088 38428 44140 38437
rect 47860 38428 47912 38480
rect 49884 38471 49936 38480
rect 49884 38437 49893 38471
rect 49893 38437 49927 38471
rect 49927 38437 49936 38471
rect 49884 38428 49936 38437
rect 49976 38428 50028 38480
rect 51172 38428 51224 38480
rect 60004 38496 60056 38548
rect 60372 38496 60424 38548
rect 37188 38224 37240 38276
rect 39212 38292 39264 38344
rect 39304 38292 39356 38344
rect 39948 38335 40000 38344
rect 39948 38301 39957 38335
rect 39957 38301 39991 38335
rect 39991 38301 40000 38335
rect 39948 38292 40000 38301
rect 41880 38292 41932 38344
rect 43720 38335 43772 38344
rect 43720 38301 43729 38335
rect 43729 38301 43763 38335
rect 43763 38301 43772 38335
rect 43720 38292 43772 38301
rect 45284 38292 45336 38344
rect 45652 38292 45704 38344
rect 47124 38335 47176 38344
rect 47124 38301 47133 38335
rect 47133 38301 47167 38335
rect 47167 38301 47176 38335
rect 47124 38292 47176 38301
rect 47768 38292 47820 38344
rect 48596 38292 48648 38344
rect 41696 38224 41748 38276
rect 41052 38156 41104 38208
rect 41972 38199 42024 38208
rect 41972 38165 41981 38199
rect 41981 38165 42015 38199
rect 42015 38165 42024 38199
rect 41972 38156 42024 38165
rect 45100 38224 45152 38276
rect 51080 38292 51132 38344
rect 43720 38156 43772 38208
rect 44732 38156 44784 38208
rect 51816 38292 51868 38344
rect 51264 38224 51316 38276
rect 51448 38156 51500 38208
rect 52276 38156 52328 38208
rect 52920 38292 52972 38344
rect 53380 38360 53432 38412
rect 54024 38428 54076 38480
rect 54484 38471 54536 38480
rect 54484 38437 54493 38471
rect 54493 38437 54527 38471
rect 54527 38437 54536 38471
rect 54484 38428 54536 38437
rect 59268 38428 59320 38480
rect 59544 38471 59596 38480
rect 59544 38437 59553 38471
rect 59553 38437 59587 38471
rect 59587 38437 59596 38471
rect 59544 38428 59596 38437
rect 53932 38360 53984 38412
rect 55220 38360 55272 38412
rect 55772 38360 55824 38412
rect 54668 38335 54720 38344
rect 54668 38301 54677 38335
rect 54677 38301 54711 38335
rect 54711 38301 54720 38335
rect 54668 38292 54720 38301
rect 56876 38335 56928 38344
rect 56876 38301 56885 38335
rect 56885 38301 56919 38335
rect 56919 38301 56928 38335
rect 56876 38292 56928 38301
rect 57152 38335 57204 38344
rect 57152 38301 57161 38335
rect 57161 38301 57195 38335
rect 57195 38301 57204 38335
rect 57152 38292 57204 38301
rect 53380 38156 53432 38208
rect 53840 38199 53892 38208
rect 53840 38165 53849 38199
rect 53849 38165 53883 38199
rect 53883 38165 53892 38199
rect 53840 38156 53892 38165
rect 57704 38292 57756 38344
rect 64236 38360 64288 38412
rect 60372 38335 60424 38344
rect 60372 38301 60381 38335
rect 60381 38301 60415 38335
rect 60415 38301 60424 38335
rect 60372 38292 60424 38301
rect 60556 38335 60608 38344
rect 60556 38301 60565 38335
rect 60565 38301 60599 38335
rect 60599 38301 60608 38335
rect 60556 38292 60608 38301
rect 57704 38156 57756 38208
rect 59176 38156 59228 38208
rect 60280 38224 60332 38276
rect 59912 38199 59964 38208
rect 59912 38165 59921 38199
rect 59921 38165 59955 38199
rect 59955 38165 59964 38199
rect 59912 38156 59964 38165
rect 60004 38156 60056 38208
rect 63132 38156 63184 38208
rect 1998 38054 2050 38106
rect 2062 38054 2114 38106
rect 2126 38054 2178 38106
rect 2190 38054 2242 38106
rect 2254 38054 2306 38106
rect 49998 38054 50050 38106
rect 50062 38054 50114 38106
rect 50126 38054 50178 38106
rect 50190 38054 50242 38106
rect 50254 38054 50306 38106
rect 7472 37995 7524 38004
rect 7472 37961 7481 37995
rect 7481 37961 7515 37995
rect 7515 37961 7524 37995
rect 7472 37952 7524 37961
rect 9312 37952 9364 38004
rect 9680 37952 9732 38004
rect 8760 37816 8812 37868
rect 11520 37952 11572 38004
rect 14372 37884 14424 37936
rect 10692 37859 10744 37868
rect 10692 37825 10701 37859
rect 10701 37825 10735 37859
rect 10735 37825 10744 37859
rect 10692 37816 10744 37825
rect 10968 37859 11020 37868
rect 10968 37825 10977 37859
rect 10977 37825 11011 37859
rect 11011 37825 11020 37859
rect 10968 37816 11020 37825
rect 13728 37816 13780 37868
rect 7564 37748 7616 37800
rect 8668 37723 8720 37732
rect 8668 37689 8677 37723
rect 8677 37689 8711 37723
rect 8711 37689 8720 37723
rect 8668 37680 8720 37689
rect 9956 37680 10008 37732
rect 10968 37612 11020 37664
rect 12256 37748 12308 37800
rect 12624 37680 12676 37732
rect 14280 37680 14332 37732
rect 14556 37859 14608 37868
rect 14556 37825 14565 37859
rect 14565 37825 14599 37859
rect 14599 37825 14608 37859
rect 14556 37816 14608 37825
rect 16488 37884 16540 37936
rect 17592 37952 17644 38004
rect 18144 37952 18196 38004
rect 18788 37952 18840 38004
rect 19340 37952 19392 38004
rect 19616 37952 19668 38004
rect 14832 37816 14884 37868
rect 15200 37859 15252 37868
rect 15200 37825 15209 37859
rect 15209 37825 15243 37859
rect 15243 37825 15252 37859
rect 15200 37816 15252 37825
rect 17776 37884 17828 37936
rect 17868 37884 17920 37936
rect 20628 37952 20680 38004
rect 20720 37952 20772 38004
rect 20996 37952 21048 38004
rect 23572 37952 23624 38004
rect 26332 37952 26384 38004
rect 26516 37952 26568 38004
rect 27804 37952 27856 38004
rect 32036 37952 32088 38004
rect 18144 37748 18196 37800
rect 18512 37791 18564 37800
rect 18512 37757 18521 37791
rect 18521 37757 18555 37791
rect 18555 37757 18564 37791
rect 18512 37748 18564 37757
rect 14096 37655 14148 37664
rect 14096 37621 14105 37655
rect 14105 37621 14139 37655
rect 14139 37621 14148 37655
rect 14096 37612 14148 37621
rect 15384 37612 15436 37664
rect 18788 37612 18840 37664
rect 19064 37655 19116 37664
rect 19064 37621 19073 37655
rect 19073 37621 19107 37655
rect 19107 37621 19116 37655
rect 19064 37612 19116 37621
rect 28264 37927 28316 37936
rect 28264 37893 28273 37927
rect 28273 37893 28307 37927
rect 28307 37893 28316 37927
rect 28264 37884 28316 37893
rect 28908 37884 28960 37936
rect 31208 37884 31260 37936
rect 33692 37952 33744 38004
rect 33968 37952 34020 38004
rect 36268 37952 36320 38004
rect 36912 37995 36964 38004
rect 36912 37961 36921 37995
rect 36921 37961 36955 37995
rect 36955 37961 36964 37995
rect 36912 37952 36964 37961
rect 37004 37952 37056 38004
rect 36452 37884 36504 37936
rect 41236 37995 41288 38004
rect 41236 37961 41245 37995
rect 41245 37961 41279 37995
rect 41279 37961 41288 37995
rect 41236 37952 41288 37961
rect 42708 37952 42760 38004
rect 43444 37952 43496 38004
rect 44548 37995 44600 38004
rect 44548 37961 44557 37995
rect 44557 37961 44591 37995
rect 44591 37961 44600 37995
rect 44548 37952 44600 37961
rect 50804 37952 50856 38004
rect 51816 37995 51868 38004
rect 51816 37961 51825 37995
rect 51825 37961 51859 37995
rect 51859 37961 51868 37995
rect 51816 37952 51868 37961
rect 26240 37816 26292 37868
rect 26792 37859 26844 37868
rect 26792 37825 26801 37859
rect 26801 37825 26835 37859
rect 26835 37825 26844 37859
rect 26792 37816 26844 37825
rect 27160 37816 27212 37868
rect 31392 37816 31444 37868
rect 31760 37816 31812 37868
rect 32312 37816 32364 37868
rect 20168 37791 20220 37800
rect 20168 37757 20177 37791
rect 20177 37757 20211 37791
rect 20211 37757 20220 37791
rect 20168 37748 20220 37757
rect 23388 37748 23440 37800
rect 28264 37748 28316 37800
rect 20812 37680 20864 37732
rect 20904 37723 20956 37732
rect 20904 37689 20913 37723
rect 20913 37689 20947 37723
rect 20947 37689 20956 37723
rect 20904 37680 20956 37689
rect 21364 37680 21416 37732
rect 19340 37612 19392 37664
rect 20260 37655 20312 37664
rect 20260 37621 20269 37655
rect 20269 37621 20303 37655
rect 20303 37621 20312 37655
rect 20260 37612 20312 37621
rect 21732 37612 21784 37664
rect 24216 37655 24268 37664
rect 24216 37621 24225 37655
rect 24225 37621 24259 37655
rect 24259 37621 24268 37655
rect 24216 37612 24268 37621
rect 24952 37723 25004 37732
rect 24952 37689 24961 37723
rect 24961 37689 24995 37723
rect 24995 37689 25004 37723
rect 24952 37680 25004 37689
rect 25044 37680 25096 37732
rect 26332 37680 26384 37732
rect 24860 37612 24912 37664
rect 26424 37655 26476 37664
rect 26424 37621 26433 37655
rect 26433 37621 26467 37655
rect 26467 37621 26476 37655
rect 26424 37612 26476 37621
rect 28080 37680 28132 37732
rect 28448 37612 28500 37664
rect 30196 37723 30248 37732
rect 30196 37689 30205 37723
rect 30205 37689 30239 37723
rect 30239 37689 30248 37723
rect 30196 37680 30248 37689
rect 32220 37680 32272 37732
rect 32404 37680 32456 37732
rect 33784 37816 33836 37868
rect 34244 37859 34296 37868
rect 34244 37825 34253 37859
rect 34253 37825 34287 37859
rect 34287 37825 34296 37859
rect 34244 37816 34296 37825
rect 34704 37816 34756 37868
rect 34980 37816 35032 37868
rect 35164 37816 35216 37868
rect 35532 37816 35584 37868
rect 33968 37748 34020 37800
rect 33876 37680 33928 37732
rect 35256 37748 35308 37800
rect 35900 37748 35952 37800
rect 37740 37748 37792 37800
rect 35164 37680 35216 37732
rect 35348 37723 35400 37732
rect 35348 37689 35357 37723
rect 35357 37689 35391 37723
rect 35391 37689 35400 37723
rect 35348 37680 35400 37689
rect 37004 37680 37056 37732
rect 39488 37816 39540 37868
rect 40776 37859 40828 37868
rect 40776 37825 40785 37859
rect 40785 37825 40819 37859
rect 40819 37825 40828 37859
rect 40776 37816 40828 37825
rect 38292 37748 38344 37800
rect 39120 37748 39172 37800
rect 40132 37748 40184 37800
rect 40500 37791 40552 37800
rect 40500 37757 40509 37791
rect 40509 37757 40543 37791
rect 40543 37757 40552 37791
rect 40500 37748 40552 37757
rect 31208 37612 31260 37664
rect 31668 37655 31720 37664
rect 31668 37621 31677 37655
rect 31677 37621 31711 37655
rect 31711 37621 31720 37655
rect 31668 37612 31720 37621
rect 32036 37612 32088 37664
rect 34704 37612 34756 37664
rect 34888 37655 34940 37664
rect 34888 37621 34897 37655
rect 34897 37621 34931 37655
rect 34931 37621 34940 37655
rect 34888 37612 34940 37621
rect 36176 37612 36228 37664
rect 37280 37612 37332 37664
rect 39304 37655 39356 37664
rect 39304 37621 39313 37655
rect 39313 37621 39347 37655
rect 39347 37621 39356 37655
rect 39304 37612 39356 37621
rect 40132 37655 40184 37664
rect 40132 37621 40141 37655
rect 40141 37621 40175 37655
rect 40175 37621 40184 37655
rect 40132 37612 40184 37621
rect 40960 37748 41012 37800
rect 42800 37816 42852 37868
rect 43352 37816 43404 37868
rect 45284 37816 45336 37868
rect 41512 37748 41564 37800
rect 41972 37748 42024 37800
rect 42708 37748 42760 37800
rect 43260 37791 43312 37800
rect 43260 37757 43269 37791
rect 43269 37757 43303 37791
rect 43303 37757 43312 37791
rect 43260 37748 43312 37757
rect 46940 37748 46992 37800
rect 48320 37816 48372 37868
rect 48412 37859 48464 37868
rect 48412 37825 48421 37859
rect 48421 37825 48455 37859
rect 48455 37825 48464 37859
rect 48412 37816 48464 37825
rect 41604 37612 41656 37664
rect 42156 37612 42208 37664
rect 45284 37680 45336 37732
rect 46020 37723 46072 37732
rect 46020 37689 46029 37723
rect 46029 37689 46063 37723
rect 46063 37689 46072 37723
rect 46020 37680 46072 37689
rect 46940 37655 46992 37664
rect 46940 37621 46949 37655
rect 46949 37621 46983 37655
rect 46983 37621 46992 37655
rect 46940 37612 46992 37621
rect 48320 37680 48372 37732
rect 49332 37791 49384 37800
rect 49332 37757 49341 37791
rect 49341 37757 49375 37791
rect 49375 37757 49384 37791
rect 49332 37748 49384 37757
rect 51356 37816 51408 37868
rect 57152 37952 57204 38004
rect 57796 37995 57848 38004
rect 57796 37961 57805 37995
rect 57805 37961 57839 37995
rect 57839 37961 57848 37995
rect 57796 37952 57848 37961
rect 55956 37884 56008 37936
rect 54668 37816 54720 37868
rect 56232 37859 56284 37868
rect 56232 37825 56241 37859
rect 56241 37825 56275 37859
rect 56275 37825 56284 37859
rect 56232 37816 56284 37825
rect 56876 37927 56928 37936
rect 56876 37893 56885 37927
rect 56885 37893 56919 37927
rect 56919 37893 56928 37927
rect 56876 37884 56928 37893
rect 58164 37859 58216 37868
rect 58164 37825 58173 37859
rect 58173 37825 58207 37859
rect 58207 37825 58216 37859
rect 58164 37816 58216 37825
rect 58256 37816 58308 37868
rect 60372 37952 60424 38004
rect 53012 37748 53064 37800
rect 55220 37748 55272 37800
rect 50344 37723 50396 37732
rect 50344 37689 50353 37723
rect 50353 37689 50387 37723
rect 50387 37689 50396 37723
rect 50344 37680 50396 37689
rect 52552 37723 52604 37732
rect 52552 37689 52561 37723
rect 52561 37689 52595 37723
rect 52595 37689 52604 37723
rect 52552 37680 52604 37689
rect 54300 37723 54352 37732
rect 54300 37689 54309 37723
rect 54309 37689 54343 37723
rect 54343 37689 54352 37723
rect 54300 37680 54352 37689
rect 56048 37748 56100 37800
rect 59268 37748 59320 37800
rect 48228 37612 48280 37664
rect 53656 37612 53708 37664
rect 56784 37680 56836 37732
rect 56876 37680 56928 37732
rect 58256 37680 58308 37732
rect 63960 37816 64012 37868
rect 60280 37791 60332 37800
rect 60280 37757 60289 37791
rect 60289 37757 60323 37791
rect 60323 37757 60332 37791
rect 60280 37748 60332 37757
rect 62488 37748 62540 37800
rect 63408 37791 63460 37800
rect 63408 37757 63417 37791
rect 63417 37757 63451 37791
rect 63451 37757 63460 37791
rect 63408 37748 63460 37757
rect 58072 37612 58124 37664
rect 59636 37655 59688 37664
rect 59636 37621 59645 37655
rect 59645 37621 59679 37655
rect 59679 37621 59688 37655
rect 59636 37612 59688 37621
rect 59820 37612 59872 37664
rect 64052 37655 64104 37664
rect 64052 37621 64061 37655
rect 64061 37621 64095 37655
rect 64095 37621 64104 37655
rect 64052 37612 64104 37621
rect 2918 37510 2970 37562
rect 2982 37510 3034 37562
rect 3046 37510 3098 37562
rect 3110 37510 3162 37562
rect 3174 37510 3226 37562
rect 50918 37510 50970 37562
rect 50982 37510 51034 37562
rect 51046 37510 51098 37562
rect 51110 37510 51162 37562
rect 51174 37510 51226 37562
rect 65258 37510 65310 37562
rect 65322 37510 65374 37562
rect 65386 37510 65438 37562
rect 65450 37510 65502 37562
rect 65514 37510 65566 37562
rect 8668 37408 8720 37460
rect 9680 37408 9732 37460
rect 10968 37451 11020 37460
rect 10968 37417 10977 37451
rect 10977 37417 11011 37451
rect 11011 37417 11020 37451
rect 10968 37408 11020 37417
rect 11336 37408 11388 37460
rect 8852 37340 8904 37392
rect 11520 37340 11572 37392
rect 12348 37340 12400 37392
rect 12624 37383 12676 37392
rect 12624 37349 12633 37383
rect 12633 37349 12667 37383
rect 12667 37349 12676 37383
rect 12624 37340 12676 37349
rect 14096 37340 14148 37392
rect 14280 37340 14332 37392
rect 15292 37451 15344 37460
rect 15292 37417 15301 37451
rect 15301 37417 15335 37451
rect 15335 37417 15344 37451
rect 15292 37408 15344 37417
rect 17684 37408 17736 37460
rect 18420 37408 18472 37460
rect 20260 37408 20312 37460
rect 21732 37451 21784 37460
rect 21732 37417 21741 37451
rect 21741 37417 21775 37451
rect 21775 37417 21784 37451
rect 21732 37408 21784 37417
rect 24952 37408 25004 37460
rect 25872 37451 25924 37460
rect 25872 37417 25881 37451
rect 25881 37417 25915 37451
rect 25915 37417 25924 37451
rect 25872 37408 25924 37417
rect 25964 37451 26016 37460
rect 25964 37417 25973 37451
rect 25973 37417 26007 37451
rect 26007 37417 26016 37451
rect 25964 37408 26016 37417
rect 26148 37408 26200 37460
rect 27436 37408 27488 37460
rect 27712 37408 27764 37460
rect 28908 37408 28960 37460
rect 30196 37408 30248 37460
rect 30748 37451 30800 37460
rect 30748 37417 30757 37451
rect 30757 37417 30791 37451
rect 30791 37417 30800 37451
rect 30748 37408 30800 37417
rect 30840 37408 30892 37460
rect 32312 37408 32364 37460
rect 32404 37451 32456 37460
rect 32404 37417 32413 37451
rect 32413 37417 32447 37451
rect 32447 37417 32456 37451
rect 32404 37408 32456 37417
rect 20720 37340 20772 37392
rect 13544 37315 13596 37324
rect 13544 37281 13553 37315
rect 13553 37281 13587 37315
rect 13587 37281 13596 37315
rect 13544 37272 13596 37281
rect 16764 37315 16816 37324
rect 16764 37281 16773 37315
rect 16773 37281 16807 37315
rect 16807 37281 16816 37315
rect 16764 37272 16816 37281
rect 18144 37272 18196 37324
rect 9588 37247 9640 37256
rect 9588 37213 9597 37247
rect 9597 37213 9631 37247
rect 9631 37213 9640 37247
rect 9588 37204 9640 37213
rect 11244 37204 11296 37256
rect 19064 37272 19116 37324
rect 23204 37272 23256 37324
rect 25044 37272 25096 37324
rect 26332 37272 26384 37324
rect 26424 37272 26476 37324
rect 30748 37272 30800 37324
rect 31668 37272 31720 37324
rect 33324 37340 33376 37392
rect 36452 37408 36504 37460
rect 36820 37408 36872 37460
rect 33508 37340 33560 37392
rect 34980 37340 35032 37392
rect 35164 37340 35216 37392
rect 36728 37383 36780 37392
rect 36728 37349 36737 37383
rect 36737 37349 36771 37383
rect 36771 37349 36780 37383
rect 36728 37340 36780 37349
rect 33600 37315 33652 37324
rect 33600 37281 33609 37315
rect 33609 37281 33643 37315
rect 33643 37281 33652 37315
rect 33600 37272 33652 37281
rect 34796 37315 34848 37324
rect 34796 37281 34805 37315
rect 34805 37281 34839 37315
rect 34839 37281 34848 37315
rect 34796 37272 34848 37281
rect 41696 37408 41748 37460
rect 42708 37408 42760 37460
rect 44916 37408 44968 37460
rect 45652 37451 45704 37460
rect 45652 37417 45661 37451
rect 45661 37417 45695 37451
rect 45695 37417 45704 37451
rect 45652 37408 45704 37417
rect 46020 37451 46072 37460
rect 46020 37417 46029 37451
rect 46029 37417 46063 37451
rect 46063 37417 46072 37451
rect 46020 37408 46072 37417
rect 47768 37451 47820 37460
rect 47768 37417 47777 37451
rect 47777 37417 47811 37451
rect 47811 37417 47820 37451
rect 47768 37408 47820 37417
rect 48228 37451 48280 37460
rect 48228 37417 48237 37451
rect 48237 37417 48271 37451
rect 48271 37417 48280 37451
rect 48228 37408 48280 37417
rect 48504 37408 48556 37460
rect 50252 37408 50304 37460
rect 50344 37408 50396 37460
rect 51264 37451 51316 37460
rect 51264 37417 51273 37451
rect 51273 37417 51307 37451
rect 51307 37417 51316 37451
rect 51264 37408 51316 37417
rect 52276 37408 52328 37460
rect 52736 37408 52788 37460
rect 53196 37451 53248 37460
rect 53196 37417 53205 37451
rect 53205 37417 53239 37451
rect 53239 37417 53248 37451
rect 53196 37408 53248 37417
rect 53564 37408 53616 37460
rect 54300 37408 54352 37460
rect 56692 37451 56744 37460
rect 56692 37417 56701 37451
rect 56701 37417 56735 37451
rect 56735 37417 56744 37451
rect 56692 37408 56744 37417
rect 58072 37408 58124 37460
rect 40132 37340 40184 37392
rect 44088 37340 44140 37392
rect 41236 37272 41288 37324
rect 41328 37272 41380 37324
rect 19248 37247 19300 37256
rect 19248 37213 19257 37247
rect 19257 37213 19291 37247
rect 19291 37213 19300 37247
rect 19248 37204 19300 37213
rect 20812 37204 20864 37256
rect 20628 37136 20680 37188
rect 25228 37136 25280 37188
rect 26516 37204 26568 37256
rect 28724 37204 28776 37256
rect 31484 37204 31536 37256
rect 27528 37136 27580 37188
rect 30288 37136 30340 37188
rect 33140 37204 33192 37256
rect 35072 37204 35124 37256
rect 35716 37204 35768 37256
rect 38476 37247 38528 37256
rect 38476 37213 38485 37247
rect 38485 37213 38519 37247
rect 38519 37213 38528 37247
rect 38476 37204 38528 37213
rect 43352 37272 43404 37324
rect 44640 37272 44692 37324
rect 44824 37315 44876 37324
rect 44824 37281 44833 37315
rect 44833 37281 44867 37315
rect 44867 37281 44876 37315
rect 44824 37272 44876 37281
rect 45100 37340 45152 37392
rect 45560 37383 45612 37392
rect 45560 37349 45569 37383
rect 45569 37349 45603 37383
rect 45603 37349 45612 37383
rect 45560 37340 45612 37349
rect 46940 37340 46992 37392
rect 49332 37340 49384 37392
rect 51816 37340 51868 37392
rect 42800 37204 42852 37256
rect 45744 37204 45796 37256
rect 47216 37247 47268 37256
rect 47216 37213 47225 37247
rect 47225 37213 47259 37247
rect 47259 37213 47268 37247
rect 47216 37204 47268 37213
rect 46756 37136 46808 37188
rect 26976 37068 27028 37120
rect 38660 37068 38712 37120
rect 41696 37111 41748 37120
rect 41696 37077 41705 37111
rect 41705 37077 41739 37111
rect 41739 37077 41748 37111
rect 41696 37068 41748 37077
rect 47124 37068 47176 37120
rect 48596 37204 48648 37256
rect 52920 37272 52972 37324
rect 56048 37315 56100 37324
rect 56048 37281 56057 37315
rect 56057 37281 56091 37315
rect 56091 37281 56100 37315
rect 56048 37272 56100 37281
rect 57152 37272 57204 37324
rect 58992 37272 59044 37324
rect 59268 37408 59320 37460
rect 59820 37340 59872 37392
rect 62488 37451 62540 37460
rect 62488 37417 62497 37451
rect 62497 37417 62531 37451
rect 62531 37417 62540 37451
rect 62488 37408 62540 37417
rect 65800 37408 65852 37460
rect 62488 37272 62540 37324
rect 64236 37315 64288 37324
rect 64236 37281 64245 37315
rect 64245 37281 64279 37315
rect 64279 37281 64288 37315
rect 64236 37272 64288 37281
rect 48688 37136 48740 37188
rect 53196 37136 53248 37188
rect 56232 37204 56284 37256
rect 56600 37247 56652 37256
rect 56600 37213 56609 37247
rect 56609 37213 56643 37247
rect 56643 37213 56652 37247
rect 56600 37204 56652 37213
rect 53748 37136 53800 37188
rect 63868 37204 63920 37256
rect 65708 37204 65760 37256
rect 54668 37068 54720 37120
rect 65432 37111 65484 37120
rect 65432 37077 65441 37111
rect 65441 37077 65475 37111
rect 65475 37077 65484 37111
rect 65432 37068 65484 37077
rect 1998 36966 2050 37018
rect 2062 36966 2114 37018
rect 2126 36966 2178 37018
rect 2190 36966 2242 37018
rect 2254 36966 2306 37018
rect 49998 36966 50050 37018
rect 50062 36966 50114 37018
rect 50126 36966 50178 37018
rect 50190 36966 50242 37018
rect 50254 36966 50306 37018
rect 64338 36966 64390 37018
rect 64402 36966 64454 37018
rect 64466 36966 64518 37018
rect 64530 36966 64582 37018
rect 64594 36966 64646 37018
rect 23480 36864 23532 36916
rect 29000 36864 29052 36916
rect 31300 36864 31352 36916
rect 35716 36864 35768 36916
rect 42248 36864 42300 36916
rect 21180 36796 21232 36848
rect 44088 36796 44140 36848
rect 47216 36864 47268 36916
rect 48596 36864 48648 36916
rect 62856 36864 62908 36916
rect 63868 36907 63920 36916
rect 63868 36873 63877 36907
rect 63877 36873 63911 36907
rect 63911 36873 63920 36907
rect 63868 36864 63920 36873
rect 22008 36728 22060 36780
rect 46756 36728 46808 36780
rect 38844 36660 38896 36712
rect 66168 36796 66220 36848
rect 60648 36728 60700 36780
rect 66536 36728 66588 36780
rect 64052 36660 64104 36712
rect 65432 36660 65484 36712
rect 24860 36592 24912 36644
rect 34428 36592 34480 36644
rect 37280 36592 37332 36644
rect 11704 36524 11756 36576
rect 8484 36456 8536 36508
rect 52552 36456 52604 36508
rect 21548 36388 21600 36440
rect 29000 36388 29052 36440
rect 30288 36320 30340 36372
rect 33048 36320 33100 36372
rect 44088 36252 44140 36304
rect 64788 36592 64840 36644
rect 64144 36524 64196 36576
rect 65156 36567 65208 36576
rect 65156 36533 65165 36567
rect 65165 36533 65199 36567
rect 65199 36533 65208 36567
rect 65156 36524 65208 36533
rect 65258 36422 65310 36474
rect 65322 36422 65374 36474
rect 65386 36422 65438 36474
rect 65450 36422 65502 36474
rect 65514 36422 65566 36474
rect 66076 36320 66128 36372
rect 25872 36184 25924 36236
rect 61568 36252 61620 36304
rect 63224 36252 63276 36304
rect 63500 36252 63552 36304
rect 64144 36295 64196 36304
rect 64144 36261 64153 36295
rect 64153 36261 64187 36295
rect 64187 36261 64196 36295
rect 64144 36252 64196 36261
rect 65800 36252 65852 36304
rect 27620 36116 27672 36168
rect 43536 36116 43588 36168
rect 63684 36184 63736 36236
rect 63776 36116 63828 36168
rect 63868 36159 63920 36168
rect 63868 36125 63877 36159
rect 63877 36125 63911 36159
rect 63911 36125 63920 36159
rect 63868 36116 63920 36125
rect 23204 36048 23256 36100
rect 38660 36048 38712 36100
rect 24676 35980 24728 36032
rect 28540 35980 28592 36032
rect 29092 35980 29144 36032
rect 62580 35980 62632 36032
rect 65708 35980 65760 36032
rect 20076 35844 20128 35896
rect 23112 35844 23164 35896
rect 23572 35844 23624 35896
rect 35808 35912 35860 35964
rect 30012 35844 30064 35896
rect 44088 35844 44140 35896
rect 64338 35878 64390 35930
rect 64402 35878 64454 35930
rect 64466 35878 64518 35930
rect 64530 35878 64582 35930
rect 64594 35878 64646 35930
rect 29000 35776 29052 35828
rect 33140 35776 33192 35828
rect 35716 35776 35768 35828
rect 40040 35776 40092 35828
rect 60556 35776 60608 35828
rect 23020 35708 23072 35760
rect 29092 35708 29144 35760
rect 31576 35708 31628 35760
rect 33600 35708 33652 35760
rect 63592 35640 63644 35692
rect 65156 35776 65208 35828
rect 63960 35708 64012 35760
rect 65156 35640 65208 35692
rect 65524 35683 65576 35692
rect 65524 35649 65533 35683
rect 65533 35649 65567 35683
rect 65567 35649 65576 35683
rect 65524 35640 65576 35649
rect 65616 35683 65668 35692
rect 65616 35649 65625 35683
rect 65625 35649 65659 35683
rect 65659 35649 65668 35683
rect 65616 35640 65668 35649
rect 61568 35572 61620 35624
rect 62488 35572 62540 35624
rect 63776 35572 63828 35624
rect 63960 35572 64012 35624
rect 8208 35504 8260 35556
rect 18052 35504 18104 35556
rect 22192 35504 22244 35556
rect 64052 35504 64104 35556
rect 65984 35504 66036 35556
rect 64144 35436 64196 35488
rect 64696 35479 64748 35488
rect 64696 35445 64705 35479
rect 64705 35445 64739 35479
rect 64739 35445 64748 35479
rect 64696 35436 64748 35445
rect 65258 35334 65310 35386
rect 65322 35334 65374 35386
rect 65386 35334 65438 35386
rect 65450 35334 65502 35386
rect 65514 35334 65566 35386
rect 62948 35232 63000 35284
rect 65616 35232 65668 35284
rect 65892 35232 65944 35284
rect 64144 35207 64196 35216
rect 64144 35173 64153 35207
rect 64153 35173 64187 35207
rect 64187 35173 64196 35207
rect 64144 35164 64196 35173
rect 65800 35164 65852 35216
rect 63868 35071 63920 35080
rect 63868 35037 63877 35071
rect 63877 35037 63911 35071
rect 63911 35037 63920 35071
rect 63868 35028 63920 35037
rect 64144 35028 64196 35080
rect 64604 35028 64656 35080
rect 65156 34892 65208 34944
rect 65616 34935 65668 34944
rect 65616 34901 65625 34935
rect 65625 34901 65659 34935
rect 65659 34901 65668 34935
rect 65616 34892 65668 34901
rect 64338 34790 64390 34842
rect 64402 34790 64454 34842
rect 64466 34790 64518 34842
rect 64530 34790 64582 34842
rect 64594 34790 64646 34842
rect 64696 34731 64748 34740
rect 64696 34697 64705 34731
rect 64705 34697 64739 34731
rect 64739 34697 64748 34731
rect 64696 34688 64748 34697
rect 62948 34552 63000 34604
rect 64788 34620 64840 34672
rect 66260 34620 66312 34672
rect 65248 34595 65300 34604
rect 65248 34561 65257 34595
rect 65257 34561 65291 34595
rect 65291 34561 65300 34595
rect 65248 34552 65300 34561
rect 65616 34484 65668 34536
rect 64052 34416 64104 34468
rect 64328 34416 64380 34468
rect 63684 34348 63736 34400
rect 64788 34348 64840 34400
rect 65258 34246 65310 34298
rect 65322 34246 65374 34298
rect 65386 34246 65438 34298
rect 65450 34246 65502 34298
rect 65514 34246 65566 34298
rect 63960 34144 64012 34196
rect 63408 34076 63460 34128
rect 64328 34076 64380 34128
rect 65616 34008 65668 34060
rect 63224 33940 63276 33992
rect 64144 33940 64196 33992
rect 63776 33804 63828 33856
rect 64972 33804 65024 33856
rect 64338 33702 64390 33754
rect 64402 33702 64454 33754
rect 64466 33702 64518 33754
rect 64530 33702 64582 33754
rect 64594 33702 64646 33754
rect 66536 33532 66588 33584
rect 65984 33507 66036 33516
rect 65984 33473 65993 33507
rect 65993 33473 66027 33507
rect 66027 33473 66036 33507
rect 65984 33464 66036 33473
rect 64328 33260 64380 33312
rect 64972 33303 65024 33312
rect 64972 33269 64981 33303
rect 64981 33269 65015 33303
rect 65015 33269 65024 33303
rect 64972 33260 65024 33269
rect 65258 33158 65310 33210
rect 65322 33158 65374 33210
rect 65386 33158 65438 33210
rect 65450 33158 65502 33210
rect 65514 33158 65566 33210
rect 65984 33056 66036 33108
rect 64236 32988 64288 33040
rect 64328 33031 64380 33040
rect 64328 32997 64337 33031
rect 64337 32997 64371 33031
rect 64371 32997 64380 33031
rect 64328 32988 64380 32997
rect 66352 32988 66404 33040
rect 64052 32963 64104 32972
rect 64052 32929 64061 32963
rect 64061 32929 64095 32963
rect 64095 32929 64104 32963
rect 64052 32920 64104 32929
rect 64338 32614 64390 32666
rect 64402 32614 64454 32666
rect 64466 32614 64518 32666
rect 64530 32614 64582 32666
rect 64594 32614 64646 32666
rect 64972 32512 65024 32564
rect 65892 32444 65944 32496
rect 65708 32376 65760 32428
rect 64696 32351 64748 32360
rect 64696 32317 64705 32351
rect 64705 32317 64739 32351
rect 64739 32317 64748 32351
rect 64696 32308 64748 32317
rect 64972 32172 65024 32224
rect 65984 32172 66036 32224
rect 65258 32070 65310 32122
rect 65322 32070 65374 32122
rect 65386 32070 65438 32122
rect 65450 32070 65502 32122
rect 65514 32070 65566 32122
rect 65800 31968 65852 32020
rect 64972 31832 65024 31884
rect 65616 31900 65668 31952
rect 65340 31832 65392 31884
rect 65892 31832 65944 31884
rect 66444 31832 66496 31884
rect 65248 31764 65300 31816
rect 64972 31696 65024 31748
rect 65708 31764 65760 31816
rect 66168 31764 66220 31816
rect 65984 31696 66036 31748
rect 64338 31526 64390 31578
rect 64402 31526 64454 31578
rect 64466 31526 64518 31578
rect 64530 31526 64582 31578
rect 64594 31526 64646 31578
rect 64052 31424 64104 31476
rect 64972 31220 65024 31272
rect 65064 31220 65116 31272
rect 65248 31220 65300 31272
rect 65258 30982 65310 31034
rect 65322 30982 65374 31034
rect 65386 30982 65438 31034
rect 65450 30982 65502 31034
rect 65514 30982 65566 31034
rect 65156 30923 65208 30932
rect 65156 30889 65165 30923
rect 65165 30889 65199 30923
rect 65199 30889 65208 30923
rect 65156 30880 65208 30889
rect 63868 30787 63920 30796
rect 63868 30753 63877 30787
rect 63877 30753 63911 30787
rect 63911 30753 63920 30787
rect 63868 30744 63920 30753
rect 64880 30744 64932 30796
rect 64880 30608 64932 30660
rect 65064 30608 65116 30660
rect 64338 30438 64390 30490
rect 64402 30438 64454 30490
rect 64466 30438 64518 30490
rect 64530 30438 64582 30490
rect 64594 30438 64646 30490
rect 65064 30200 65116 30252
rect 64328 30107 64380 30116
rect 64328 30073 64337 30107
rect 64337 30073 64371 30107
rect 64371 30073 64380 30107
rect 64328 30064 64380 30073
rect 66444 30064 66496 30116
rect 65984 29996 66036 30048
rect 62948 29928 63000 29980
rect 63132 29928 63184 29980
rect 65258 29894 65310 29946
rect 65322 29894 65374 29946
rect 65386 29894 65438 29946
rect 65450 29894 65502 29946
rect 65514 29894 65566 29946
rect 64328 29792 64380 29844
rect 65708 29835 65760 29844
rect 65708 29801 65717 29835
rect 65717 29801 65751 29835
rect 65751 29801 65760 29835
rect 65708 29792 65760 29801
rect 65800 29835 65852 29844
rect 65800 29801 65809 29835
rect 65809 29801 65843 29835
rect 65843 29801 65852 29835
rect 65800 29792 65852 29801
rect 65064 29724 65116 29776
rect 65156 29656 65208 29708
rect 66536 29588 66588 29640
rect 64696 29452 64748 29504
rect 64338 29350 64390 29402
rect 64402 29350 64454 29402
rect 64466 29350 64518 29402
rect 64530 29350 64582 29402
rect 64594 29350 64646 29402
rect 65616 29248 65668 29300
rect 64052 29155 64104 29164
rect 64052 29121 64061 29155
rect 64061 29121 64095 29155
rect 64095 29121 64104 29155
rect 64052 29112 64104 29121
rect 64696 29112 64748 29164
rect 65800 28976 65852 29028
rect 66444 28976 66496 29028
rect 65258 28806 65310 28858
rect 65322 28806 65374 28858
rect 65386 28806 65438 28858
rect 65450 28806 65502 28858
rect 65514 28806 65566 28858
rect 63316 28704 63368 28756
rect 65156 28747 65208 28756
rect 65156 28713 65165 28747
rect 65165 28713 65199 28747
rect 65199 28713 65208 28747
rect 65156 28704 65208 28713
rect 65064 28636 65116 28688
rect 65984 28704 66036 28756
rect 65616 28568 65668 28620
rect 64880 28432 64932 28484
rect 65156 28432 65208 28484
rect 64338 28262 64390 28314
rect 64402 28262 64454 28314
rect 64466 28262 64518 28314
rect 64530 28262 64582 28314
rect 64594 28262 64646 28314
rect 63316 28160 63368 28212
rect 65258 27718 65310 27770
rect 65322 27718 65374 27770
rect 65386 27718 65438 27770
rect 65450 27718 65502 27770
rect 65514 27718 65566 27770
rect 65616 27616 65668 27668
rect 64880 27480 64932 27532
rect 65156 27412 65208 27464
rect 65708 27412 65760 27464
rect 65064 27276 65116 27328
rect 64338 27174 64390 27226
rect 64402 27174 64454 27226
rect 64466 27174 64518 27226
rect 64530 27174 64582 27226
rect 64594 27174 64646 27226
rect 64696 26936 64748 26988
rect 65800 26868 65852 26920
rect 65984 26868 66036 26920
rect 64604 26800 64656 26852
rect 65800 26775 65852 26784
rect 65800 26741 65809 26775
rect 65809 26741 65843 26775
rect 65843 26741 65852 26775
rect 65800 26732 65852 26741
rect 65258 26630 65310 26682
rect 65322 26630 65374 26682
rect 65386 26630 65438 26682
rect 65450 26630 65502 26682
rect 65514 26630 65566 26682
rect 64604 26571 64656 26580
rect 64604 26537 64613 26571
rect 64613 26537 64647 26571
rect 64647 26537 64656 26571
rect 64604 26528 64656 26537
rect 65064 26571 65116 26580
rect 65064 26537 65073 26571
rect 65073 26537 65107 26571
rect 65107 26537 65116 26571
rect 65064 26528 65116 26537
rect 65524 26528 65576 26580
rect 65984 26528 66036 26580
rect 65800 26392 65852 26444
rect 65984 26435 66036 26444
rect 65984 26401 65993 26435
rect 65993 26401 66027 26435
rect 66027 26401 66036 26435
rect 65984 26392 66036 26401
rect 65156 26324 65208 26376
rect 66536 26324 66588 26376
rect 64880 26256 64932 26308
rect 65800 26256 65852 26308
rect 63868 26188 63920 26240
rect 64052 26188 64104 26240
rect 64338 26086 64390 26138
rect 64402 26086 64454 26138
rect 64466 26086 64518 26138
rect 64530 26086 64582 26138
rect 64594 26086 64646 26138
rect 65258 25542 65310 25594
rect 65322 25542 65374 25594
rect 65386 25542 65438 25594
rect 65450 25542 65502 25594
rect 65514 25542 65566 25594
rect 63960 25347 64012 25356
rect 63960 25313 63969 25347
rect 63969 25313 64003 25347
rect 64003 25313 64012 25347
rect 63960 25304 64012 25313
rect 65064 25279 65116 25288
rect 65064 25245 65073 25279
rect 65073 25245 65107 25279
rect 65107 25245 65116 25279
rect 65064 25236 65116 25245
rect 65156 25279 65208 25288
rect 65156 25245 65165 25279
rect 65165 25245 65199 25279
rect 65199 25245 65208 25279
rect 65156 25236 65208 25245
rect 65800 25236 65852 25288
rect 64236 25100 64288 25152
rect 64338 24998 64390 25050
rect 64402 24998 64454 25050
rect 64466 24998 64518 25050
rect 64530 24998 64582 25050
rect 64594 24998 64646 25050
rect 63224 24828 63276 24880
rect 63592 24828 63644 24880
rect 64972 24692 65024 24744
rect 63960 24556 64012 24608
rect 65258 24454 65310 24506
rect 65322 24454 65374 24506
rect 65386 24454 65438 24506
rect 65450 24454 65502 24506
rect 65514 24454 65566 24506
rect 64696 24352 64748 24404
rect 64052 24284 64104 24336
rect 64338 23910 64390 23962
rect 64402 23910 64454 23962
rect 64466 23910 64518 23962
rect 64530 23910 64582 23962
rect 64594 23910 64646 23962
rect 63960 23604 64012 23656
rect 64236 23536 64288 23588
rect 65616 23536 65668 23588
rect 63040 23468 63092 23520
rect 63868 23468 63920 23520
rect 65800 23511 65852 23520
rect 65800 23477 65809 23511
rect 65809 23477 65843 23511
rect 65843 23477 65852 23511
rect 65800 23468 65852 23477
rect 65258 23366 65310 23418
rect 65322 23366 65374 23418
rect 65386 23366 65438 23418
rect 65450 23366 65502 23418
rect 65514 23366 65566 23418
rect 65064 23264 65116 23316
rect 65984 23196 66036 23248
rect 64880 23171 64932 23180
rect 64880 23137 64889 23171
rect 64889 23137 64923 23171
rect 64923 23137 64932 23171
rect 64880 23128 64932 23137
rect 65892 23128 65944 23180
rect 65708 23060 65760 23112
rect 64338 22822 64390 22874
rect 64402 22822 64454 22874
rect 64466 22822 64518 22874
rect 64530 22822 64582 22874
rect 64594 22822 64646 22874
rect 64880 22720 64932 22772
rect 64052 22516 64104 22568
rect 64696 22516 64748 22568
rect 64144 22448 64196 22500
rect 64880 22448 64932 22500
rect 65892 22448 65944 22500
rect 65258 22278 65310 22330
rect 65322 22278 65374 22330
rect 65386 22278 65438 22330
rect 65450 22278 65502 22330
rect 65514 22278 65566 22330
rect 66260 22176 66312 22228
rect 65892 22108 65944 22160
rect 63960 22040 64012 22092
rect 64696 21972 64748 22024
rect 64338 21734 64390 21786
rect 64402 21734 64454 21786
rect 64466 21734 64518 21786
rect 64530 21734 64582 21786
rect 64594 21734 64646 21786
rect 65708 21428 65760 21480
rect 66260 21428 66312 21480
rect 63316 21360 63368 21412
rect 63868 21360 63920 21412
rect 65616 21360 65668 21412
rect 65156 21292 65208 21344
rect 65258 21190 65310 21242
rect 65322 21190 65374 21242
rect 65386 21190 65438 21242
rect 65450 21190 65502 21242
rect 65514 21190 65566 21242
rect 64696 21088 64748 21140
rect 65156 21088 65208 21140
rect 65064 20927 65116 20936
rect 65064 20893 65073 20927
rect 65073 20893 65107 20927
rect 65107 20893 65116 20927
rect 65064 20884 65116 20893
rect 65616 20884 65668 20936
rect 64338 20646 64390 20698
rect 64402 20646 64454 20698
rect 64466 20646 64518 20698
rect 64530 20646 64582 20698
rect 64594 20646 64646 20698
rect 64972 20408 65024 20460
rect 65800 20340 65852 20392
rect 64144 20272 64196 20324
rect 66168 20272 66220 20324
rect 64880 20204 64932 20256
rect 65800 20204 65852 20256
rect 65258 20102 65310 20154
rect 65322 20102 65374 20154
rect 65386 20102 65438 20154
rect 65450 20102 65502 20154
rect 65514 20102 65566 20154
rect 65892 19932 65944 19984
rect 66168 19932 66220 19984
rect 64052 19839 64104 19848
rect 64052 19805 64061 19839
rect 64061 19805 64095 19839
rect 64095 19805 64104 19839
rect 64052 19796 64104 19805
rect 64696 19796 64748 19848
rect 65892 19660 65944 19712
rect 64338 19558 64390 19610
rect 64402 19558 64454 19610
rect 64466 19558 64518 19610
rect 64530 19558 64582 19610
rect 64594 19558 64646 19610
rect 64696 19456 64748 19508
rect 65616 19320 65668 19372
rect 64880 19252 64932 19304
rect 65892 19252 65944 19304
rect 65258 19014 65310 19066
rect 65322 19014 65374 19066
rect 65386 19014 65438 19066
rect 65450 19014 65502 19066
rect 65514 19014 65566 19066
rect 65064 18751 65116 18760
rect 65064 18717 65073 18751
rect 65073 18717 65107 18751
rect 65107 18717 65116 18751
rect 65064 18708 65116 18717
rect 65616 18708 65668 18760
rect 65984 18751 66036 18760
rect 65984 18717 65993 18751
rect 65993 18717 66027 18751
rect 66027 18717 66036 18751
rect 65984 18708 66036 18717
rect 64696 18572 64748 18624
rect 64338 18470 64390 18522
rect 64402 18470 64454 18522
rect 64466 18470 64518 18522
rect 64530 18470 64582 18522
rect 64594 18470 64646 18522
rect 63040 18368 63092 18420
rect 66076 18368 66128 18420
rect 64696 18232 64748 18284
rect 64052 18207 64104 18216
rect 64052 18173 64061 18207
rect 64061 18173 64095 18207
rect 64095 18173 64104 18207
rect 64052 18164 64104 18173
rect 66168 18096 66220 18148
rect 64972 18028 65024 18080
rect 65984 18028 66036 18080
rect 65258 17926 65310 17978
rect 65322 17926 65374 17978
rect 65386 17926 65438 17978
rect 65450 17926 65502 17978
rect 65514 17926 65566 17978
rect 64972 17824 65024 17876
rect 65064 17824 65116 17876
rect 65708 17867 65760 17876
rect 65708 17833 65717 17867
rect 65717 17833 65751 17867
rect 65751 17833 65760 17867
rect 65708 17824 65760 17833
rect 64696 17756 64748 17808
rect 65984 17688 66036 17740
rect 64880 17620 64932 17672
rect 65156 17552 65208 17604
rect 64338 17382 64390 17434
rect 64402 17382 64454 17434
rect 64466 17382 64518 17434
rect 64530 17382 64582 17434
rect 64594 17382 64646 17434
rect 64696 17280 64748 17332
rect 65258 16838 65310 16890
rect 65322 16838 65374 16890
rect 65386 16838 65438 16890
rect 65450 16838 65502 16890
rect 65514 16838 65566 16890
rect 62948 16668 63000 16720
rect 66076 16668 66128 16720
rect 63316 16600 63368 16652
rect 65800 16600 65852 16652
rect 65064 16575 65116 16584
rect 65064 16541 65073 16575
rect 65073 16541 65107 16575
rect 65107 16541 65116 16575
rect 65064 16532 65116 16541
rect 63500 16396 63552 16448
rect 64696 16396 64748 16448
rect 64338 16294 64390 16346
rect 64402 16294 64454 16346
rect 64466 16294 64518 16346
rect 64530 16294 64582 16346
rect 64594 16294 64646 16346
rect 65800 16235 65852 16244
rect 65800 16201 65809 16235
rect 65809 16201 65843 16235
rect 65843 16201 65852 16235
rect 65800 16192 65852 16201
rect 63960 16056 64012 16108
rect 64696 16056 64748 16108
rect 66168 15920 66220 15972
rect 65258 15750 65310 15802
rect 65322 15750 65374 15802
rect 65386 15750 65438 15802
rect 65450 15750 65502 15802
rect 65514 15750 65566 15802
rect 64788 15648 64840 15700
rect 65064 15648 65116 15700
rect 65892 15580 65944 15632
rect 64880 15444 64932 15496
rect 65156 15444 65208 15496
rect 64338 15206 64390 15258
rect 64402 15206 64454 15258
rect 64466 15206 64518 15258
rect 64530 15206 64582 15258
rect 64594 15206 64646 15258
rect 64788 15104 64840 15156
rect 65258 14662 65310 14714
rect 65322 14662 65374 14714
rect 65386 14662 65438 14714
rect 65450 14662 65502 14714
rect 65514 14662 65566 14714
rect 64338 14118 64390 14170
rect 64402 14118 64454 14170
rect 64466 14118 64518 14170
rect 64530 14118 64582 14170
rect 64594 14118 64646 14170
rect 65258 13574 65310 13626
rect 65322 13574 65374 13626
rect 65386 13574 65438 13626
rect 65450 13574 65502 13626
rect 65514 13574 65566 13626
rect 64338 13030 64390 13082
rect 64402 13030 64454 13082
rect 64466 13030 64518 13082
rect 64530 13030 64582 13082
rect 64594 13030 64646 13082
rect 63960 12792 64012 12844
rect 65064 12792 65116 12844
rect 66076 12835 66128 12844
rect 66076 12801 66085 12835
rect 66085 12801 66119 12835
rect 66119 12801 66128 12835
rect 66076 12792 66128 12801
rect 64788 12656 64840 12708
rect 66444 12588 66496 12640
rect 65258 12486 65310 12538
rect 65322 12486 65374 12538
rect 65386 12486 65438 12538
rect 65450 12486 65502 12538
rect 65514 12486 65566 12538
rect 65984 12384 66036 12436
rect 66168 12316 66220 12368
rect 63868 12180 63920 12232
rect 64696 12180 64748 12232
rect 64338 11942 64390 11994
rect 64402 11942 64454 11994
rect 64466 11942 64518 11994
rect 64530 11942 64582 11994
rect 64594 11942 64646 11994
rect 64696 11840 64748 11892
rect 65064 11840 65116 11892
rect 65616 11704 65668 11756
rect 62948 11636 63000 11688
rect 64144 11636 64196 11688
rect 66260 11636 66312 11688
rect 66076 11568 66128 11620
rect 64880 11543 64932 11552
rect 64880 11509 64889 11543
rect 64889 11509 64923 11543
rect 64923 11509 64932 11543
rect 64880 11500 64932 11509
rect 65892 11500 65944 11552
rect 65258 11398 65310 11450
rect 65322 11398 65374 11450
rect 65386 11398 65438 11450
rect 65450 11398 65502 11450
rect 65514 11398 65566 11450
rect 64880 11296 64932 11348
rect 65984 11203 66036 11212
rect 65984 11169 65993 11203
rect 65993 11169 66027 11203
rect 66027 11169 66036 11203
rect 65984 11160 66036 11169
rect 64338 10854 64390 10906
rect 64402 10854 64454 10906
rect 64466 10854 64518 10906
rect 64530 10854 64582 10906
rect 64594 10854 64646 10906
rect 65616 10684 65668 10736
rect 65156 10659 65208 10668
rect 65156 10625 65165 10659
rect 65165 10625 65199 10659
rect 65199 10625 65208 10659
rect 65156 10616 65208 10625
rect 65800 10548 65852 10600
rect 64972 10455 65024 10464
rect 64972 10421 64981 10455
rect 64981 10421 65015 10455
rect 65015 10421 65024 10455
rect 64972 10412 65024 10421
rect 65258 10310 65310 10362
rect 65322 10310 65374 10362
rect 65386 10310 65438 10362
rect 65450 10310 65502 10362
rect 65514 10310 65566 10362
rect 66168 10140 66220 10192
rect 63868 10004 63920 10056
rect 64696 10004 64748 10056
rect 64972 9868 65024 9920
rect 64338 9766 64390 9818
rect 64402 9766 64454 9818
rect 64466 9766 64518 9818
rect 64530 9766 64582 9818
rect 64594 9766 64646 9818
rect 63224 9596 63276 9648
rect 63960 9596 64012 9648
rect 65156 9571 65208 9580
rect 65156 9537 65191 9571
rect 65191 9537 65208 9571
rect 65156 9528 65208 9537
rect 64880 9460 64932 9512
rect 64972 9460 65024 9512
rect 65064 9392 65116 9444
rect 64972 9367 65024 9376
rect 64972 9333 64981 9367
rect 64981 9333 65015 9367
rect 65015 9333 65024 9367
rect 64972 9324 65024 9333
rect 65156 9324 65208 9376
rect 65258 9222 65310 9274
rect 65322 9222 65374 9274
rect 65386 9222 65438 9274
rect 65450 9222 65502 9274
rect 65514 9222 65566 9274
rect 64696 9120 64748 9172
rect 65064 9120 65116 9172
rect 64972 8984 65024 9036
rect 65984 8984 66036 9036
rect 63500 8916 63552 8968
rect 64236 8916 64288 8968
rect 65064 8959 65116 8968
rect 65064 8925 65073 8959
rect 65073 8925 65107 8959
rect 65107 8925 65116 8959
rect 65064 8916 65116 8925
rect 65248 8959 65300 8968
rect 65248 8925 65257 8959
rect 65257 8925 65291 8959
rect 65291 8925 65300 8959
rect 65248 8916 65300 8925
rect 65708 8916 65760 8968
rect 64338 8678 64390 8730
rect 64402 8678 64454 8730
rect 64466 8678 64518 8730
rect 64530 8678 64582 8730
rect 64594 8678 64646 8730
rect 65248 8483 65300 8492
rect 65248 8449 65257 8483
rect 65257 8449 65291 8483
rect 65291 8449 65300 8483
rect 65248 8440 65300 8449
rect 65616 8372 65668 8424
rect 65800 8372 65852 8424
rect 64604 8279 64656 8288
rect 64604 8245 64613 8279
rect 64613 8245 64647 8279
rect 64647 8245 64656 8279
rect 64604 8236 64656 8245
rect 65258 8134 65310 8186
rect 65322 8134 65374 8186
rect 65386 8134 65438 8186
rect 65450 8134 65502 8186
rect 65514 8134 65566 8186
rect 64604 7964 64656 8016
rect 66168 7964 66220 8016
rect 64052 7939 64104 7948
rect 64052 7905 64061 7939
rect 64061 7905 64095 7939
rect 64095 7905 64104 7939
rect 64052 7896 64104 7905
rect 65800 7735 65852 7744
rect 65800 7701 65809 7735
rect 65809 7701 65843 7735
rect 65843 7701 65852 7735
rect 65800 7692 65852 7701
rect 64338 7590 64390 7642
rect 64402 7590 64454 7642
rect 64466 7590 64518 7642
rect 64530 7590 64582 7642
rect 64594 7590 64646 7642
rect 65064 7488 65116 7540
rect 64880 7420 64932 7472
rect 65800 7352 65852 7404
rect 64512 7284 64564 7336
rect 65984 7327 66036 7336
rect 65984 7293 65993 7327
rect 65993 7293 66027 7327
rect 66027 7293 66036 7327
rect 65984 7284 66036 7293
rect 65616 7148 65668 7200
rect 65258 7046 65310 7098
rect 65322 7046 65374 7098
rect 65386 7046 65438 7098
rect 65450 7046 65502 7098
rect 65514 7046 65566 7098
rect 65616 6944 65668 6996
rect 62856 6808 62908 6860
rect 63592 6808 63644 6860
rect 64512 6851 64564 6860
rect 64512 6817 64521 6851
rect 64521 6817 64555 6851
rect 64555 6817 64564 6851
rect 64512 6808 64564 6817
rect 64604 6808 64656 6860
rect 65156 6808 65208 6860
rect 64972 6740 65024 6792
rect 65616 6740 65668 6792
rect 64788 6604 64840 6656
rect 64338 6502 64390 6554
rect 64402 6502 64454 6554
rect 64466 6502 64518 6554
rect 64530 6502 64582 6554
rect 64594 6502 64646 6554
rect 66260 6400 66312 6452
rect 64144 6332 64196 6384
rect 64512 6332 64564 6384
rect 64972 6264 65024 6316
rect 63960 6196 64012 6248
rect 64512 6196 64564 6248
rect 65984 6196 66036 6248
rect 64880 6128 64932 6180
rect 64328 6060 64380 6112
rect 65258 5958 65310 6010
rect 65322 5958 65374 6010
rect 65386 5958 65438 6010
rect 65450 5958 65502 6010
rect 65514 5958 65566 6010
rect 63592 5856 63644 5908
rect 64144 5856 64196 5908
rect 64328 5899 64380 5908
rect 64328 5865 64337 5899
rect 64337 5865 64371 5899
rect 64371 5865 64380 5899
rect 64328 5856 64380 5865
rect 64512 5856 64564 5908
rect 63592 5720 63644 5772
rect 64328 5652 64380 5704
rect 63960 5516 64012 5568
rect 64338 5414 64390 5466
rect 64402 5414 64454 5466
rect 64466 5414 64518 5466
rect 64530 5414 64582 5466
rect 64594 5414 64646 5466
rect 65984 5312 66036 5364
rect 64052 5219 64104 5228
rect 64052 5185 64061 5219
rect 64061 5185 64095 5219
rect 64095 5185 64104 5219
rect 64052 5176 64104 5185
rect 64788 5176 64840 5228
rect 65708 5040 65760 5092
rect 66168 5040 66220 5092
rect 65258 4870 65310 4922
rect 65322 4870 65374 4922
rect 65386 4870 65438 4922
rect 65450 4870 65502 4922
rect 65514 4870 65566 4922
rect 64880 4768 64932 4820
rect 65156 4768 65208 4820
rect 65708 4700 65760 4752
rect 63868 4675 63920 4684
rect 63868 4641 63877 4675
rect 63877 4641 63911 4675
rect 63911 4641 63920 4675
rect 63868 4632 63920 4641
rect 64696 4564 64748 4616
rect 64338 4326 64390 4378
rect 64402 4326 64454 4378
rect 64466 4326 64518 4378
rect 64530 4326 64582 4378
rect 64594 4326 64646 4378
rect 63960 4224 64012 4276
rect 64052 3952 64104 4004
rect 66444 3952 66496 4004
rect 64144 3884 64196 3936
rect 65258 3782 65310 3834
rect 65322 3782 65374 3834
rect 65386 3782 65438 3834
rect 65450 3782 65502 3834
rect 65514 3782 65566 3834
rect 64144 3723 64196 3732
rect 64144 3689 64153 3723
rect 64153 3689 64187 3723
rect 64187 3689 64196 3723
rect 64144 3680 64196 3689
rect 63500 3612 63552 3664
rect 63868 3612 63920 3664
rect 65064 3587 65116 3596
rect 65064 3553 65073 3587
rect 65073 3553 65107 3587
rect 65107 3553 65116 3587
rect 65064 3544 65116 3553
rect 65616 3476 65668 3528
rect 64972 3408 65024 3460
rect 64696 3383 64748 3392
rect 64696 3349 64705 3383
rect 64705 3349 64739 3383
rect 64739 3349 64748 3383
rect 64696 3340 64748 3349
rect 64338 3238 64390 3290
rect 64402 3238 64454 3290
rect 64466 3238 64518 3290
rect 64530 3238 64582 3290
rect 64594 3238 64646 3290
rect 63868 3179 63920 3188
rect 63868 3145 63877 3179
rect 63877 3145 63911 3179
rect 63911 3145 63920 3179
rect 63868 3136 63920 3145
rect 64052 3043 64104 3052
rect 64052 3009 64061 3043
rect 64061 3009 64095 3043
rect 64095 3009 64104 3043
rect 64052 3000 64104 3009
rect 64236 2864 64288 2916
rect 65708 2864 65760 2916
rect 65800 2839 65852 2848
rect 65800 2805 65809 2839
rect 65809 2805 65843 2839
rect 65843 2805 65852 2839
rect 65800 2796 65852 2805
rect 65258 2694 65310 2746
rect 65322 2694 65374 2746
rect 65386 2694 65438 2746
rect 65450 2694 65502 2746
rect 65514 2694 65566 2746
rect 63592 2592 63644 2644
rect 64972 2592 65024 2644
rect 66076 2592 66128 2644
rect 64144 2456 64196 2508
rect 65156 2456 65208 2508
rect 64328 2388 64380 2440
rect 64696 2388 64748 2440
rect 64788 2295 64840 2304
rect 64788 2261 64797 2295
rect 64797 2261 64831 2295
rect 64831 2261 64840 2295
rect 64788 2252 64840 2261
rect 64338 2150 64390 2202
rect 64402 2150 64454 2202
rect 64466 2150 64518 2202
rect 64530 2150 64582 2202
rect 64594 2150 64646 2202
rect 65064 2048 65116 2100
rect 48964 1980 49016 2032
rect 63040 1980 63092 2032
rect 65892 1980 65944 2032
rect 49608 1912 49660 1964
rect 62488 1912 62540 1964
rect 64696 1955 64748 1964
rect 64696 1921 64705 1955
rect 64705 1921 64739 1955
rect 64739 1921 64748 1955
rect 64696 1912 64748 1921
rect 65800 1912 65852 1964
rect 49700 1844 49752 1896
rect 63776 1844 63828 1896
rect 65156 1844 65208 1896
rect 64696 1776 64748 1828
rect 64972 1819 65024 1828
rect 64972 1785 64981 1819
rect 64981 1785 65015 1819
rect 65015 1785 65024 1819
rect 64972 1776 65024 1785
rect 65258 1606 65310 1658
rect 65322 1606 65374 1658
rect 65386 1606 65438 1658
rect 65450 1606 65502 1658
rect 65514 1606 65566 1658
rect 64696 1547 64748 1556
rect 64696 1513 64705 1547
rect 64705 1513 64739 1547
rect 64739 1513 64748 1547
rect 64696 1504 64748 1513
rect 64788 1504 64840 1556
rect 64236 1368 64288 1420
rect 65156 1411 65208 1420
rect 65156 1377 65165 1411
rect 65165 1377 65199 1411
rect 65199 1377 65208 1411
rect 65156 1368 65208 1377
rect 65616 1300 65668 1352
rect 64338 1062 64390 1114
rect 64402 1062 64454 1114
rect 64466 1062 64518 1114
rect 64530 1062 64582 1114
rect 64594 1062 64646 1114
rect 65156 960 65208 1012
rect 65800 824 65852 876
rect 65258 518 65310 570
rect 65322 518 65374 570
rect 65386 518 65438 570
rect 65450 518 65502 570
rect 65514 518 65566 570
<< metal2 >>
rect 34610 45112 34666 45121
rect 34610 45047 34666 45056
rect 21272 45008 21324 45014
rect 21272 44950 21324 44956
rect 11702 44840 11758 44849
rect 11702 44775 11758 44784
rect 13818 44840 13874 44849
rect 13818 44775 13874 44784
rect 15108 44804 15160 44810
rect 11150 44704 11206 44713
rect 1998 44636 2306 44645
rect 11150 44639 11206 44648
rect 1998 44634 2004 44636
rect 2060 44634 2084 44636
rect 2140 44634 2164 44636
rect 2220 44634 2244 44636
rect 2300 44634 2306 44636
rect 2060 44582 2062 44634
rect 2242 44582 2244 44634
rect 1998 44580 2004 44582
rect 2060 44580 2084 44582
rect 2140 44580 2164 44582
rect 2220 44580 2244 44582
rect 2300 44580 2306 44582
rect 1998 44571 2306 44580
rect 6182 44568 6238 44577
rect 6182 44503 6184 44512
rect 6236 44503 6238 44512
rect 6734 44568 6790 44577
rect 6734 44503 6736 44512
rect 6184 44474 6236 44480
rect 6788 44503 6790 44512
rect 7286 44568 7342 44577
rect 7286 44503 7288 44512
rect 6736 44474 6788 44480
rect 7340 44503 7342 44512
rect 7838 44568 7894 44577
rect 7838 44503 7840 44512
rect 7288 44474 7340 44480
rect 7892 44503 7894 44512
rect 8390 44568 8446 44577
rect 8390 44503 8392 44512
rect 7840 44474 7892 44480
rect 8444 44503 8446 44512
rect 8942 44568 8998 44577
rect 8942 44503 8944 44512
rect 8392 44474 8444 44480
rect 8996 44503 8998 44512
rect 9494 44568 9550 44577
rect 9494 44503 9496 44512
rect 8944 44474 8996 44480
rect 9548 44503 9550 44512
rect 10046 44568 10102 44577
rect 10046 44503 10048 44512
rect 9496 44474 9548 44480
rect 10100 44503 10102 44512
rect 10506 44568 10562 44577
rect 10506 44503 10508 44512
rect 10048 44474 10100 44480
rect 10560 44503 10562 44512
rect 10782 44568 10838 44577
rect 11164 44538 11192 44639
rect 11426 44568 11482 44577
rect 10782 44503 10784 44512
rect 10508 44474 10560 44480
rect 10836 44503 10838 44512
rect 11152 44532 11204 44538
rect 10784 44474 10836 44480
rect 11716 44538 11744 44775
rect 12530 44568 12586 44577
rect 11426 44503 11428 44512
rect 11152 44474 11204 44480
rect 11480 44503 11482 44512
rect 11704 44532 11756 44538
rect 11428 44474 11480 44480
rect 12530 44503 12532 44512
rect 11704 44474 11756 44480
rect 12584 44503 12586 44512
rect 12532 44474 12584 44480
rect 13832 44470 13860 44775
rect 15108 44746 15160 44752
rect 14556 44736 14608 44742
rect 14370 44704 14426 44713
rect 14556 44678 14608 44684
rect 14370 44639 14426 44648
rect 13820 44464 13872 44470
rect 13820 44406 13872 44412
rect 14384 44334 14412 44639
rect 14568 44334 14596 44678
rect 15120 44334 15148 44746
rect 15198 44568 15254 44577
rect 20074 44568 20130 44577
rect 15198 44503 15200 44512
rect 15252 44503 15254 44512
rect 18420 44532 18472 44538
rect 15200 44474 15252 44480
rect 20074 44503 20076 44512
rect 18420 44474 18472 44480
rect 20128 44503 20130 44512
rect 20076 44474 20128 44480
rect 16488 44464 16540 44470
rect 16488 44406 16540 44412
rect 14372 44328 14424 44334
rect 14372 44270 14424 44276
rect 14556 44328 14608 44334
rect 14556 44270 14608 44276
rect 15108 44328 15160 44334
rect 15108 44270 15160 44276
rect 15384 44328 15436 44334
rect 15384 44270 15436 44276
rect 14096 44260 14148 44266
rect 14096 44202 14148 44208
rect 11612 44192 11664 44198
rect 11612 44134 11664 44140
rect 13728 44192 13780 44198
rect 13728 44134 13780 44140
rect 2918 44092 3226 44101
rect 2918 44090 2924 44092
rect 2980 44090 3004 44092
rect 3060 44090 3084 44092
rect 3140 44090 3164 44092
rect 3220 44090 3226 44092
rect 2980 44038 2982 44090
rect 3162 44038 3164 44090
rect 2918 44036 2924 44038
rect 2980 44036 3004 44038
rect 3060 44036 3084 44038
rect 3140 44036 3164 44038
rect 3220 44036 3226 44038
rect 2918 44027 3226 44036
rect 11624 43790 11652 44134
rect 13740 44010 13768 44134
rect 13648 43982 13768 44010
rect 12532 43920 12584 43926
rect 12532 43862 12584 43868
rect 12806 43888 12862 43897
rect 11612 43784 11664 43790
rect 11612 43726 11664 43732
rect 11704 43784 11756 43790
rect 11704 43726 11756 43732
rect 11060 43648 11112 43654
rect 11060 43590 11112 43596
rect 1998 43548 2306 43557
rect 1998 43546 2004 43548
rect 2060 43546 2084 43548
rect 2140 43546 2164 43548
rect 2220 43546 2244 43548
rect 2300 43546 2306 43548
rect 2060 43494 2062 43546
rect 2242 43494 2244 43546
rect 1998 43492 2004 43494
rect 2060 43492 2084 43494
rect 2140 43492 2164 43494
rect 2220 43492 2244 43494
rect 2300 43492 2306 43494
rect 1998 43483 2306 43492
rect 10692 43240 10744 43246
rect 10692 43182 10744 43188
rect 2918 43004 3226 43013
rect 2918 43002 2924 43004
rect 2980 43002 3004 43004
rect 3060 43002 3084 43004
rect 3140 43002 3164 43004
rect 3220 43002 3226 43004
rect 2980 42950 2982 43002
rect 3162 42950 3164 43002
rect 2918 42948 2924 42950
rect 2980 42948 3004 42950
rect 3060 42948 3084 42950
rect 3140 42948 3164 42950
rect 3220 42948 3226 42950
rect 2918 42939 3226 42948
rect 9496 42696 9548 42702
rect 9496 42638 9548 42644
rect 8944 42560 8996 42566
rect 8944 42502 8996 42508
rect 1998 42460 2306 42469
rect 1998 42458 2004 42460
rect 2060 42458 2084 42460
rect 2140 42458 2164 42460
rect 2220 42458 2244 42460
rect 2300 42458 2306 42460
rect 2060 42406 2062 42458
rect 2242 42406 2244 42458
rect 1998 42404 2004 42406
rect 2060 42404 2084 42406
rect 2140 42404 2164 42406
rect 2220 42404 2244 42406
rect 2300 42404 2306 42406
rect 1998 42395 2306 42404
rect 8392 42220 8444 42226
rect 8392 42162 8444 42168
rect 2918 41916 3226 41925
rect 2918 41914 2924 41916
rect 2980 41914 3004 41916
rect 3060 41914 3084 41916
rect 3140 41914 3164 41916
rect 3220 41914 3226 41916
rect 2980 41862 2982 41914
rect 3162 41862 3164 41914
rect 2918 41860 2924 41862
rect 2980 41860 3004 41862
rect 3060 41860 3084 41862
rect 3140 41860 3164 41862
rect 3220 41860 3226 41862
rect 2918 41851 3226 41860
rect 8300 41744 8352 41750
rect 8404 41732 8432 42162
rect 8576 42016 8628 42022
rect 8576 41958 8628 41964
rect 8352 41704 8432 41732
rect 8300 41686 8352 41692
rect 8024 41608 8076 41614
rect 8024 41550 8076 41556
rect 1998 41372 2306 41381
rect 1998 41370 2004 41372
rect 2060 41370 2084 41372
rect 2140 41370 2164 41372
rect 2220 41370 2244 41372
rect 2300 41370 2306 41372
rect 2060 41318 2062 41370
rect 2242 41318 2244 41370
rect 1998 41316 2004 41318
rect 2060 41316 2084 41318
rect 2140 41316 2164 41318
rect 2220 41316 2244 41318
rect 2300 41316 2306 41318
rect 1998 41307 2306 41316
rect 7748 40928 7800 40934
rect 7748 40870 7800 40876
rect 2918 40828 3226 40837
rect 2918 40826 2924 40828
rect 2980 40826 3004 40828
rect 3060 40826 3084 40828
rect 3140 40826 3164 40828
rect 3220 40826 3226 40828
rect 2980 40774 2982 40826
rect 3162 40774 3164 40826
rect 2918 40772 2924 40774
rect 2980 40772 3004 40774
rect 3060 40772 3084 40774
rect 3140 40772 3164 40774
rect 3220 40772 3226 40774
rect 2918 40763 3226 40772
rect 7760 40390 7788 40870
rect 8036 40730 8064 41550
rect 8404 41138 8432 41704
rect 8300 41132 8352 41138
rect 8300 41074 8352 41080
rect 8392 41132 8444 41138
rect 8392 41074 8444 41080
rect 8024 40724 8076 40730
rect 8024 40666 8076 40672
rect 8312 40594 8340 41074
rect 8300 40588 8352 40594
rect 8300 40530 8352 40536
rect 7748 40384 7800 40390
rect 7748 40326 7800 40332
rect 1998 40284 2306 40293
rect 1998 40282 2004 40284
rect 2060 40282 2084 40284
rect 2140 40282 2164 40284
rect 2220 40282 2244 40284
rect 2300 40282 2306 40284
rect 2060 40230 2062 40282
rect 2242 40230 2244 40282
rect 1998 40228 2004 40230
rect 2060 40228 2084 40230
rect 2140 40228 2164 40230
rect 2220 40228 2244 40230
rect 2300 40228 2306 40230
rect 1998 40219 2306 40228
rect 7656 39976 7708 39982
rect 7656 39918 7708 39924
rect 2918 39740 3226 39749
rect 2918 39738 2924 39740
rect 2980 39738 3004 39740
rect 3060 39738 3084 39740
rect 3140 39738 3164 39740
rect 3220 39738 3226 39740
rect 2980 39686 2982 39738
rect 3162 39686 3164 39738
rect 2918 39684 2924 39686
rect 2980 39684 3004 39686
rect 3060 39684 3084 39686
rect 3140 39684 3164 39686
rect 3220 39684 3226 39686
rect 2918 39675 3226 39684
rect 7668 39438 7696 39918
rect 7656 39432 7708 39438
rect 7656 39374 7708 39380
rect 1998 39196 2306 39205
rect 1998 39194 2004 39196
rect 2060 39194 2084 39196
rect 2140 39194 2164 39196
rect 2220 39194 2244 39196
rect 2300 39194 2306 39196
rect 2060 39142 2062 39194
rect 2242 39142 2244 39194
rect 1998 39140 2004 39142
rect 2060 39140 2084 39142
rect 2140 39140 2164 39142
rect 2220 39140 2244 39142
rect 2300 39140 2306 39142
rect 1998 39131 2306 39140
rect 7564 38752 7616 38758
rect 7564 38694 7616 38700
rect 2918 38652 3226 38661
rect 2918 38650 2924 38652
rect 2980 38650 3004 38652
rect 3060 38650 3084 38652
rect 3140 38650 3164 38652
rect 3220 38650 3226 38652
rect 2980 38598 2982 38650
rect 3162 38598 3164 38650
rect 2918 38596 2924 38598
rect 2980 38596 3004 38598
rect 3060 38596 3084 38598
rect 3140 38596 3164 38598
rect 3220 38596 3226 38598
rect 2918 38587 3226 38596
rect 7472 38344 7524 38350
rect 7472 38286 7524 38292
rect 1998 38108 2306 38117
rect 1998 38106 2004 38108
rect 2060 38106 2084 38108
rect 2140 38106 2164 38108
rect 2220 38106 2244 38108
rect 2300 38106 2306 38108
rect 2060 38054 2062 38106
rect 2242 38054 2244 38106
rect 1998 38052 2004 38054
rect 2060 38052 2084 38054
rect 2140 38052 2164 38054
rect 2220 38052 2244 38054
rect 2300 38052 2306 38054
rect 1998 38043 2306 38052
rect 7484 38010 7512 38286
rect 7472 38004 7524 38010
rect 7472 37946 7524 37952
rect 7576 37806 7604 38694
rect 8404 38554 8432 41074
rect 8588 41002 8616 41958
rect 8576 40996 8628 41002
rect 8576 40938 8628 40944
rect 8956 40730 8984 42502
rect 9508 41818 9536 42638
rect 9680 42152 9732 42158
rect 9680 42094 9732 42100
rect 9496 41812 9548 41818
rect 9496 41754 9548 41760
rect 9588 41676 9640 41682
rect 9588 41618 9640 41624
rect 9036 41540 9088 41546
rect 9036 41482 9088 41488
rect 8944 40724 8996 40730
rect 8944 40666 8996 40672
rect 9048 40662 9076 41482
rect 9036 40656 9088 40662
rect 9036 40598 9088 40604
rect 8576 40520 8628 40526
rect 8576 40462 8628 40468
rect 8760 40520 8812 40526
rect 8760 40462 8812 40468
rect 8588 40118 8616 40462
rect 8772 40186 8800 40462
rect 8760 40180 8812 40186
rect 8760 40122 8812 40128
rect 8576 40112 8628 40118
rect 8576 40054 8628 40060
rect 8576 39568 8628 39574
rect 8576 39510 8628 39516
rect 8588 39098 8616 39510
rect 8576 39092 8628 39098
rect 8576 39034 8628 39040
rect 8772 38962 8800 40122
rect 9312 40044 9364 40050
rect 9312 39986 9364 39992
rect 8852 39840 8904 39846
rect 8852 39782 8904 39788
rect 9128 39840 9180 39846
rect 9128 39782 9180 39788
rect 8864 39574 8892 39782
rect 8852 39568 8904 39574
rect 8852 39510 8904 39516
rect 8852 39296 8904 39302
rect 8852 39238 8904 39244
rect 8760 38956 8812 38962
rect 8760 38898 8812 38904
rect 8668 38820 8720 38826
rect 8668 38762 8720 38768
rect 8680 38554 8708 38762
rect 8392 38548 8444 38554
rect 8392 38490 8444 38496
rect 8668 38548 8720 38554
rect 8668 38490 8720 38496
rect 8772 37874 8800 38898
rect 8864 38826 8892 39238
rect 8852 38820 8904 38826
rect 8852 38762 8904 38768
rect 9140 38554 9168 39782
rect 8852 38548 8904 38554
rect 8852 38490 8904 38496
rect 9128 38548 9180 38554
rect 9128 38490 9180 38496
rect 8760 37868 8812 37874
rect 8760 37810 8812 37816
rect 7564 37800 7616 37806
rect 7564 37742 7616 37748
rect 8668 37732 8720 37738
rect 8668 37674 8720 37680
rect 2918 37564 3226 37573
rect 2918 37562 2924 37564
rect 2980 37562 3004 37564
rect 3060 37562 3084 37564
rect 3140 37562 3164 37564
rect 3220 37562 3226 37564
rect 2980 37510 2982 37562
rect 3162 37510 3164 37562
rect 2918 37508 2924 37510
rect 2980 37508 3004 37510
rect 3060 37508 3084 37510
rect 3140 37508 3164 37510
rect 3220 37508 3226 37510
rect 2918 37499 3226 37508
rect 8680 37466 8708 37674
rect 8668 37460 8720 37466
rect 8668 37402 8720 37408
rect 8864 37398 8892 38490
rect 9324 38282 9352 39986
rect 9496 39568 9548 39574
rect 9496 39510 9548 39516
rect 9508 38554 9536 39510
rect 9600 39370 9628 41618
rect 9692 41274 9720 42094
rect 10324 41744 10376 41750
rect 10324 41686 10376 41692
rect 10232 41608 10284 41614
rect 10232 41550 10284 41556
rect 9680 41268 9732 41274
rect 9680 41210 9732 41216
rect 10244 41206 10272 41550
rect 10232 41200 10284 41206
rect 10232 41142 10284 41148
rect 10336 41002 10364 41686
rect 10324 40996 10376 41002
rect 10324 40938 10376 40944
rect 10232 40928 10284 40934
rect 10232 40870 10284 40876
rect 10244 40050 10272 40870
rect 10336 40662 10364 40938
rect 10324 40656 10376 40662
rect 10324 40598 10376 40604
rect 10416 40520 10468 40526
rect 10416 40462 10468 40468
rect 10232 40044 10284 40050
rect 10232 39986 10284 39992
rect 10428 39370 10456 40462
rect 10704 40458 10732 43182
rect 11072 42022 11100 43590
rect 11244 43172 11296 43178
rect 11244 43114 11296 43120
rect 11256 42906 11284 43114
rect 11244 42900 11296 42906
rect 11244 42842 11296 42848
rect 11520 42220 11572 42226
rect 11520 42162 11572 42168
rect 11060 42016 11112 42022
rect 11060 41958 11112 41964
rect 10784 41676 10836 41682
rect 10784 41618 10836 41624
rect 10796 40594 10824 41618
rect 11532 41614 11560 42162
rect 11520 41608 11572 41614
rect 11520 41550 11572 41556
rect 11336 40928 11388 40934
rect 11336 40870 11388 40876
rect 11348 40730 11376 40870
rect 11336 40724 11388 40730
rect 11336 40666 11388 40672
rect 10968 40656 11020 40662
rect 10968 40598 11020 40604
rect 10784 40588 10836 40594
rect 10784 40530 10836 40536
rect 10692 40452 10744 40458
rect 10692 40394 10744 40400
rect 10704 40202 10732 40394
rect 10520 40186 10732 40202
rect 10508 40180 10732 40186
rect 10560 40174 10732 40180
rect 10508 40122 10560 40128
rect 9588 39364 9640 39370
rect 9588 39306 9640 39312
rect 10416 39364 10468 39370
rect 10416 39306 10468 39312
rect 9496 38548 9548 38554
rect 9496 38490 9548 38496
rect 9312 38276 9364 38282
rect 9312 38218 9364 38224
rect 9324 38010 9352 38218
rect 9312 38004 9364 38010
rect 9312 37946 9364 37952
rect 8852 37392 8904 37398
rect 8852 37334 8904 37340
rect 9600 37262 9628 39306
rect 9956 38412 10008 38418
rect 9956 38354 10008 38360
rect 9680 38344 9732 38350
rect 9680 38286 9732 38292
rect 9692 38010 9720 38286
rect 9680 38004 9732 38010
rect 9680 37946 9732 37952
rect 9692 37466 9720 37946
rect 9968 37738 9996 38354
rect 10704 37874 10732 40174
rect 10980 40050 11008 40598
rect 11244 40520 11296 40526
rect 11244 40462 11296 40468
rect 10968 40044 11020 40050
rect 10968 39986 11020 39992
rect 10980 38826 11008 39986
rect 10876 38820 10928 38826
rect 10876 38762 10928 38768
rect 10968 38820 11020 38826
rect 10968 38762 11020 38768
rect 10888 38554 10916 38762
rect 11256 38554 11284 40462
rect 11348 40050 11376 40666
rect 11336 40044 11388 40050
rect 11336 39986 11388 39992
rect 11426 39672 11482 39681
rect 11426 39607 11482 39616
rect 11440 39574 11468 39607
rect 11428 39568 11480 39574
rect 11428 39510 11480 39516
rect 11440 39098 11468 39510
rect 11428 39092 11480 39098
rect 11428 39034 11480 39040
rect 11532 38962 11560 41550
rect 11624 41138 11652 43726
rect 11716 42906 11744 43726
rect 12256 43716 12308 43722
rect 12256 43658 12308 43664
rect 11704 42900 11756 42906
rect 11704 42842 11756 42848
rect 11716 42362 11744 42842
rect 11704 42356 11756 42362
rect 11704 42298 11756 42304
rect 12268 42090 12296 43658
rect 12544 42362 12572 43862
rect 12806 43823 12808 43832
rect 12860 43823 12862 43832
rect 12808 43794 12860 43800
rect 13648 43738 13676 43982
rect 13728 43920 13780 43926
rect 13728 43862 13780 43868
rect 13556 43710 13676 43738
rect 12624 43648 12676 43654
rect 12624 43590 12676 43596
rect 12636 42702 12664 43590
rect 12716 43104 12768 43110
rect 12716 43046 12768 43052
rect 12992 43104 13044 43110
rect 12992 43046 13044 43052
rect 12728 42770 12756 43046
rect 12716 42764 12768 42770
rect 12716 42706 12768 42712
rect 12624 42696 12676 42702
rect 12624 42638 12676 42644
rect 12532 42356 12584 42362
rect 12532 42298 12584 42304
rect 12256 42084 12308 42090
rect 12256 42026 12308 42032
rect 11796 41608 11848 41614
rect 11796 41550 11848 41556
rect 11808 41274 11836 41550
rect 11796 41268 11848 41274
rect 11796 41210 11848 41216
rect 12072 41268 12124 41274
rect 12072 41210 12124 41216
rect 11612 41132 11664 41138
rect 11612 41074 11664 41080
rect 11704 40588 11756 40594
rect 11704 40530 11756 40536
rect 11716 39506 11744 40530
rect 12084 40526 12112 41210
rect 12072 40520 12124 40526
rect 12072 40462 12124 40468
rect 11704 39500 11756 39506
rect 11704 39442 11756 39448
rect 11520 38956 11572 38962
rect 11520 38898 11572 38904
rect 10876 38548 10928 38554
rect 10876 38490 10928 38496
rect 11244 38548 11296 38554
rect 11244 38490 11296 38496
rect 11256 38418 11284 38490
rect 11244 38412 11296 38418
rect 11244 38354 11296 38360
rect 10968 38208 11020 38214
rect 10968 38150 11020 38156
rect 10980 37874 11008 38150
rect 10692 37868 10744 37874
rect 10692 37810 10744 37816
rect 10968 37868 11020 37874
rect 10968 37810 11020 37816
rect 9956 37732 10008 37738
rect 9956 37674 10008 37680
rect 10968 37664 11020 37670
rect 10968 37606 11020 37612
rect 10980 37466 11008 37606
rect 9680 37460 9732 37466
rect 9680 37402 9732 37408
rect 10968 37460 11020 37466
rect 10968 37402 11020 37408
rect 11256 37262 11284 38354
rect 11336 38344 11388 38350
rect 11336 38286 11388 38292
rect 11348 37466 11376 38286
rect 11520 38004 11572 38010
rect 11520 37946 11572 37952
rect 11336 37460 11388 37466
rect 11336 37402 11388 37408
rect 11532 37398 11560 37946
rect 11520 37392 11572 37398
rect 11520 37334 11572 37340
rect 9588 37256 9640 37262
rect 9588 37198 9640 37204
rect 11244 37256 11296 37262
rect 11244 37198 11296 37204
rect 1998 37020 2306 37029
rect 1998 37018 2004 37020
rect 2060 37018 2084 37020
rect 2140 37018 2164 37020
rect 2220 37018 2244 37020
rect 2300 37018 2306 37020
rect 2060 36966 2062 37018
rect 2242 36966 2244 37018
rect 1998 36964 2004 36966
rect 2060 36964 2084 36966
rect 2140 36964 2164 36966
rect 2220 36964 2244 36966
rect 2300 36964 2306 36966
rect 1998 36955 2306 36964
rect 11716 36582 11744 39442
rect 12268 37806 12296 42026
rect 12440 42016 12492 42022
rect 12492 41976 12572 42004
rect 12440 41958 12492 41964
rect 12440 41472 12492 41478
rect 12440 41414 12492 41420
rect 12452 41070 12480 41414
rect 12440 41064 12492 41070
rect 12440 41006 12492 41012
rect 12440 40928 12492 40934
rect 12440 40870 12492 40876
rect 12452 40662 12480 40870
rect 12544 40662 12572 41976
rect 12636 41206 12664 42638
rect 12728 42090 12756 42706
rect 12808 42696 12860 42702
rect 12808 42638 12860 42644
rect 12716 42084 12768 42090
rect 12716 42026 12768 42032
rect 12624 41200 12676 41206
rect 12624 41142 12676 41148
rect 12440 40656 12492 40662
rect 12440 40598 12492 40604
rect 12532 40656 12584 40662
rect 12532 40598 12584 40604
rect 12544 40118 12572 40598
rect 12532 40112 12584 40118
rect 12532 40054 12584 40060
rect 12544 39658 12572 40054
rect 12452 39630 12572 39658
rect 12820 39642 12848 42638
rect 13004 42226 13032 43046
rect 13556 42566 13584 43710
rect 13636 43648 13688 43654
rect 13636 43590 13688 43596
rect 13648 43314 13676 43590
rect 13636 43308 13688 43314
rect 13636 43250 13688 43256
rect 13740 43110 13768 43862
rect 13820 43716 13872 43722
rect 13820 43658 13872 43664
rect 13832 43178 13860 43658
rect 13820 43172 13872 43178
rect 13820 43114 13872 43120
rect 13728 43104 13780 43110
rect 13728 43046 13780 43052
rect 13832 42838 13860 43114
rect 13820 42832 13872 42838
rect 13820 42774 13872 42780
rect 13176 42560 13228 42566
rect 13176 42502 13228 42508
rect 13544 42560 13596 42566
rect 13544 42502 13596 42508
rect 13188 42226 13216 42502
rect 12992 42220 13044 42226
rect 12992 42162 13044 42168
rect 13176 42220 13228 42226
rect 13176 42162 13228 42168
rect 12992 41608 13044 41614
rect 12992 41550 13044 41556
rect 12900 41132 12952 41138
rect 12900 41074 12952 41080
rect 12808 39636 12860 39642
rect 12452 39574 12480 39630
rect 12808 39578 12860 39584
rect 12440 39568 12492 39574
rect 12912 39522 12940 41074
rect 13004 41070 13032 41550
rect 13188 41414 13216 42162
rect 13728 42152 13780 42158
rect 13728 42094 13780 42100
rect 13636 42084 13688 42090
rect 13636 42026 13688 42032
rect 13188 41386 13308 41414
rect 13280 41274 13308 41386
rect 13268 41268 13320 41274
rect 13268 41210 13320 41216
rect 13280 41138 13308 41210
rect 13268 41132 13320 41138
rect 13268 41074 13320 41080
rect 12992 41064 13044 41070
rect 12992 41006 13044 41012
rect 12992 39976 13044 39982
rect 13648 39953 13676 42026
rect 13740 41206 13768 42094
rect 13832 41750 13860 42774
rect 14108 42650 14136 44202
rect 14740 44192 14792 44198
rect 14740 44134 14792 44140
rect 14648 43988 14700 43994
rect 14648 43930 14700 43936
rect 14464 43648 14516 43654
rect 14464 43590 14516 43596
rect 14476 42702 14504 43590
rect 14660 42906 14688 43930
rect 14752 43772 14780 44134
rect 15200 43920 15252 43926
rect 15200 43862 15252 43868
rect 14924 43784 14976 43790
rect 14752 43744 14924 43772
rect 14924 43726 14976 43732
rect 14648 42900 14700 42906
rect 14648 42842 14700 42848
rect 14464 42696 14516 42702
rect 14108 42622 14228 42650
rect 14464 42638 14516 42644
rect 13820 41744 13872 41750
rect 13820 41686 13872 41692
rect 13832 41414 13860 41686
rect 13832 41386 14136 41414
rect 13728 41200 13780 41206
rect 13728 41142 13780 41148
rect 13740 40050 13768 41142
rect 13820 41064 13872 41070
rect 13820 41006 13872 41012
rect 14002 41032 14058 41041
rect 13832 40526 13860 41006
rect 14002 40967 14004 40976
rect 14056 40967 14058 40976
rect 14004 40938 14056 40944
rect 13912 40928 13964 40934
rect 13912 40870 13964 40876
rect 13924 40526 13952 40870
rect 14016 40730 14044 40938
rect 14004 40724 14056 40730
rect 14004 40666 14056 40672
rect 13820 40520 13872 40526
rect 13820 40462 13872 40468
rect 13912 40520 13964 40526
rect 13912 40462 13964 40468
rect 13728 40044 13780 40050
rect 13728 39986 13780 39992
rect 12992 39918 13044 39924
rect 13634 39944 13690 39953
rect 12440 39510 12492 39516
rect 12820 39494 12940 39522
rect 12820 38962 12848 39494
rect 13004 39302 13032 39918
rect 13634 39879 13690 39888
rect 13084 39840 13136 39846
rect 13084 39782 13136 39788
rect 13096 39438 13124 39782
rect 13544 39568 13596 39574
rect 13544 39510 13596 39516
rect 13084 39432 13136 39438
rect 13084 39374 13136 39380
rect 12992 39296 13044 39302
rect 12992 39238 13044 39244
rect 12808 38956 12860 38962
rect 12808 38898 12860 38904
rect 12348 38752 12400 38758
rect 12348 38694 12400 38700
rect 12360 38418 12388 38694
rect 12348 38412 12400 38418
rect 12348 38354 12400 38360
rect 12820 38350 12848 38898
rect 13004 38894 13032 39238
rect 12992 38888 13044 38894
rect 12992 38830 13044 38836
rect 13452 38820 13504 38826
rect 13556 38808 13584 39510
rect 13504 38780 13584 38808
rect 13452 38762 13504 38768
rect 12808 38344 12860 38350
rect 12808 38286 12860 38292
rect 12624 38276 12676 38282
rect 12624 38218 12676 38224
rect 12256 37800 12308 37806
rect 12256 37742 12308 37748
rect 12636 37738 12664 38218
rect 12624 37732 12676 37738
rect 12624 37674 12676 37680
rect 12636 37505 12664 37674
rect 12622 37496 12678 37505
rect 12622 37431 12678 37440
rect 12636 37398 12664 37431
rect 12348 37392 12400 37398
rect 12348 37334 12400 37340
rect 12624 37392 12676 37398
rect 12624 37334 12676 37340
rect 12360 36689 12388 37334
rect 13556 37330 13584 38780
rect 13648 38554 13676 39879
rect 13832 38962 13860 40462
rect 13912 39908 13964 39914
rect 13912 39850 13964 39856
rect 13924 39506 13952 39850
rect 13912 39500 13964 39506
rect 13912 39442 13964 39448
rect 13820 38956 13872 38962
rect 13820 38898 13872 38904
rect 14108 38826 14136 41386
rect 14200 39846 14228 42622
rect 14372 42016 14424 42022
rect 14372 41958 14424 41964
rect 14384 41818 14412 41958
rect 14372 41812 14424 41818
rect 14372 41754 14424 41760
rect 14936 41414 14964 43726
rect 15212 42906 15240 43862
rect 15396 43450 15424 44270
rect 15936 44192 15988 44198
rect 15936 44134 15988 44140
rect 15948 43994 15976 44134
rect 15936 43988 15988 43994
rect 15936 43930 15988 43936
rect 16210 43888 16266 43897
rect 16210 43823 16212 43832
rect 16264 43823 16266 43832
rect 16212 43794 16264 43800
rect 15936 43648 15988 43654
rect 15936 43590 15988 43596
rect 15384 43444 15436 43450
rect 15384 43386 15436 43392
rect 15384 43240 15436 43246
rect 15384 43182 15436 43188
rect 15200 42900 15252 42906
rect 15200 42842 15252 42848
rect 15396 42362 15424 43182
rect 15948 43178 15976 43590
rect 15936 43172 15988 43178
rect 15936 43114 15988 43120
rect 15568 43104 15620 43110
rect 15568 43046 15620 43052
rect 15580 42838 15608 43046
rect 16500 42838 16528 44406
rect 17224 44396 17276 44402
rect 17224 44338 17276 44344
rect 16856 44192 16908 44198
rect 16856 44134 16908 44140
rect 16868 42906 16896 44134
rect 17236 43976 17264 44338
rect 17776 44328 17828 44334
rect 17776 44270 17828 44276
rect 17592 44260 17644 44266
rect 17592 44202 17644 44208
rect 17684 44260 17736 44266
rect 17684 44202 17736 44208
rect 17408 43988 17460 43994
rect 17236 43948 17408 43976
rect 17132 43648 17184 43654
rect 17132 43590 17184 43596
rect 16856 42900 16908 42906
rect 16856 42842 16908 42848
rect 17144 42838 17172 43590
rect 15568 42832 15620 42838
rect 15568 42774 15620 42780
rect 16488 42832 16540 42838
rect 16488 42774 16540 42780
rect 17132 42832 17184 42838
rect 17132 42774 17184 42780
rect 15384 42356 15436 42362
rect 15384 42298 15436 42304
rect 15580 42265 15608 42774
rect 15844 42764 15896 42770
rect 15844 42706 15896 42712
rect 15566 42256 15622 42265
rect 15566 42191 15622 42200
rect 15476 42016 15528 42022
rect 15476 41958 15528 41964
rect 15384 41472 15436 41478
rect 15384 41414 15436 41420
rect 14384 41386 14964 41414
rect 14188 39840 14240 39846
rect 14188 39782 14240 39788
rect 14384 39438 14412 41386
rect 15016 41064 15068 41070
rect 15016 41006 15068 41012
rect 14556 40928 14608 40934
rect 14556 40870 14608 40876
rect 14568 40594 14596 40870
rect 15028 40662 15056 41006
rect 15200 40996 15252 41002
rect 15200 40938 15252 40944
rect 15212 40730 15240 40938
rect 15200 40724 15252 40730
rect 15200 40666 15252 40672
rect 15016 40656 15068 40662
rect 15016 40598 15068 40604
rect 14556 40588 14608 40594
rect 14556 40530 14608 40536
rect 15292 40520 15344 40526
rect 15292 40462 15344 40468
rect 14464 39500 14516 39506
rect 14464 39442 14516 39448
rect 14372 39432 14424 39438
rect 14372 39374 14424 39380
rect 14096 38820 14148 38826
rect 14096 38762 14148 38768
rect 13636 38548 13688 38554
rect 13636 38490 13688 38496
rect 13728 38344 13780 38350
rect 13728 38286 13780 38292
rect 13740 37874 13768 38286
rect 14384 38214 14412 39374
rect 14476 38554 14504 39442
rect 15304 39438 15332 40462
rect 15396 40186 15424 41414
rect 15488 40730 15516 41958
rect 15568 41608 15620 41614
rect 15568 41550 15620 41556
rect 15660 41608 15712 41614
rect 15660 41550 15712 41556
rect 15476 40724 15528 40730
rect 15476 40666 15528 40672
rect 15580 40610 15608 41550
rect 15488 40582 15608 40610
rect 15384 40180 15436 40186
rect 15384 40122 15436 40128
rect 15488 40118 15516 40582
rect 15672 40526 15700 41550
rect 15856 41274 15884 42706
rect 16028 42628 16080 42634
rect 16028 42570 16080 42576
rect 16040 42362 16068 42570
rect 16304 42560 16356 42566
rect 16304 42502 16356 42508
rect 16396 42560 16448 42566
rect 16396 42502 16448 42508
rect 16316 42362 16344 42502
rect 16028 42356 16080 42362
rect 16028 42298 16080 42304
rect 16304 42356 16356 42362
rect 16304 42298 16356 42304
rect 16408 42226 16436 42502
rect 16396 42220 16448 42226
rect 16396 42162 16448 42168
rect 16500 41614 16528 42774
rect 17144 42702 17172 42774
rect 16672 42696 16724 42702
rect 16672 42638 16724 42644
rect 16948 42696 17000 42702
rect 16948 42638 17000 42644
rect 17132 42696 17184 42702
rect 17132 42638 17184 42644
rect 16684 42226 16712 42638
rect 16960 42362 16988 42638
rect 16948 42356 17000 42362
rect 16948 42298 17000 42304
rect 16672 42220 16724 42226
rect 16672 42162 16724 42168
rect 17236 42022 17264 43948
rect 17408 43930 17460 43936
rect 17604 43790 17632 44202
rect 17592 43784 17644 43790
rect 17592 43726 17644 43732
rect 17498 43480 17554 43489
rect 17498 43415 17500 43424
rect 17552 43415 17554 43424
rect 17500 43386 17552 43392
rect 17696 43178 17724 44202
rect 17788 43994 17816 44270
rect 18144 44192 18196 44198
rect 18144 44134 18196 44140
rect 17776 43988 17828 43994
rect 17776 43930 17828 43936
rect 17868 43784 17920 43790
rect 17868 43726 17920 43732
rect 17684 43172 17736 43178
rect 17684 43114 17736 43120
rect 17314 42936 17370 42945
rect 17696 42906 17724 43114
rect 17776 43104 17828 43110
rect 17776 43046 17828 43052
rect 17314 42871 17370 42880
rect 17684 42900 17736 42906
rect 17328 42770 17356 42871
rect 17684 42842 17736 42848
rect 17316 42764 17368 42770
rect 17316 42706 17368 42712
rect 17592 42764 17644 42770
rect 17592 42706 17644 42712
rect 17604 42566 17632 42706
rect 17592 42560 17644 42566
rect 17592 42502 17644 42508
rect 17696 42158 17724 42842
rect 17788 42838 17816 43046
rect 17776 42832 17828 42838
rect 17776 42774 17828 42780
rect 17880 42362 17908 43726
rect 18052 43376 18104 43382
rect 18052 43318 18104 43324
rect 17958 42392 18014 42401
rect 17868 42356 17920 42362
rect 17958 42327 18014 42336
rect 17868 42298 17920 42304
rect 17684 42152 17736 42158
rect 17684 42094 17736 42100
rect 17040 42016 17092 42022
rect 17040 41958 17092 41964
rect 17224 42016 17276 42022
rect 17224 41958 17276 41964
rect 17592 42016 17644 42022
rect 17592 41958 17644 41964
rect 17052 41750 17080 41958
rect 17236 41750 17264 41958
rect 16764 41744 16816 41750
rect 16764 41686 16816 41692
rect 17040 41744 17092 41750
rect 17040 41686 17092 41692
rect 17224 41744 17276 41750
rect 17224 41686 17276 41692
rect 16488 41608 16540 41614
rect 16488 41550 16540 41556
rect 16776 41274 16804 41686
rect 17132 41676 17184 41682
rect 17132 41618 17184 41624
rect 16856 41608 16908 41614
rect 16856 41550 16908 41556
rect 15844 41268 15896 41274
rect 15844 41210 15896 41216
rect 16488 41268 16540 41274
rect 16764 41268 16816 41274
rect 16540 41228 16620 41256
rect 16488 41210 16540 41216
rect 15752 40996 15804 41002
rect 15752 40938 15804 40944
rect 15660 40520 15712 40526
rect 15660 40462 15712 40468
rect 15764 40390 15792 40938
rect 15856 40594 15884 41210
rect 15844 40588 15896 40594
rect 15844 40530 15896 40536
rect 15936 40520 15988 40526
rect 15936 40462 15988 40468
rect 16488 40520 16540 40526
rect 16488 40462 16540 40468
rect 15568 40384 15620 40390
rect 15568 40326 15620 40332
rect 15752 40384 15804 40390
rect 15752 40326 15804 40332
rect 15476 40112 15528 40118
rect 15476 40054 15528 40060
rect 15476 39976 15528 39982
rect 15476 39918 15528 39924
rect 15488 39574 15516 39918
rect 15580 39574 15608 40326
rect 15764 39914 15792 40326
rect 15752 39908 15804 39914
rect 15752 39850 15804 39856
rect 15476 39568 15528 39574
rect 15476 39510 15528 39516
rect 15568 39568 15620 39574
rect 15568 39510 15620 39516
rect 15292 39432 15344 39438
rect 15292 39374 15344 39380
rect 15200 39024 15252 39030
rect 15200 38966 15252 38972
rect 14832 38956 14884 38962
rect 14832 38898 14884 38904
rect 14464 38548 14516 38554
rect 14464 38490 14516 38496
rect 14556 38276 14608 38282
rect 14556 38218 14608 38224
rect 14372 38208 14424 38214
rect 14372 38150 14424 38156
rect 14384 37942 14412 38150
rect 14372 37936 14424 37942
rect 14372 37878 14424 37884
rect 14568 37874 14596 38218
rect 14844 37874 14872 38898
rect 15212 38486 15240 38966
rect 15292 38888 15344 38894
rect 15292 38830 15344 38836
rect 15200 38480 15252 38486
rect 15200 38422 15252 38428
rect 15304 38418 15332 38830
rect 15384 38752 15436 38758
rect 15384 38694 15436 38700
rect 15292 38412 15344 38418
rect 15292 38354 15344 38360
rect 15200 38208 15252 38214
rect 15200 38150 15252 38156
rect 15212 37874 15240 38150
rect 13728 37868 13780 37874
rect 13728 37810 13780 37816
rect 14556 37868 14608 37874
rect 14556 37810 14608 37816
rect 14832 37868 14884 37874
rect 14832 37810 14884 37816
rect 15200 37868 15252 37874
rect 15200 37810 15252 37816
rect 14280 37732 14332 37738
rect 14280 37674 14332 37680
rect 14096 37664 14148 37670
rect 14096 37606 14148 37612
rect 14108 37398 14136 37606
rect 14292 37398 14320 37674
rect 15304 37466 15332 38354
rect 15396 37670 15424 38694
rect 15488 38486 15516 39510
rect 15948 39370 15976 40462
rect 16500 40050 16528 40462
rect 16488 40044 16540 40050
rect 16488 39986 16540 39992
rect 15936 39364 15988 39370
rect 15936 39306 15988 39312
rect 16396 39024 16448 39030
rect 16396 38966 16448 38972
rect 16210 38856 16266 38865
rect 16210 38791 16266 38800
rect 15476 38480 15528 38486
rect 15476 38422 15528 38428
rect 15384 37664 15436 37670
rect 15384 37606 15436 37612
rect 15292 37460 15344 37466
rect 15292 37402 15344 37408
rect 14096 37392 14148 37398
rect 14096 37334 14148 37340
rect 14280 37392 14332 37398
rect 14280 37334 14332 37340
rect 13544 37324 13596 37330
rect 13544 37266 13596 37272
rect 16224 36961 16252 38791
rect 16408 38350 16436 38966
rect 16488 38548 16540 38554
rect 16488 38490 16540 38496
rect 16500 38418 16528 38490
rect 16488 38412 16540 38418
rect 16488 38354 16540 38360
rect 16396 38344 16448 38350
rect 16396 38286 16448 38292
rect 16210 36952 16266 36961
rect 16210 36887 16266 36896
rect 16408 36689 16436 38286
rect 16500 37942 16528 38354
rect 16488 37936 16540 37942
rect 16592 37913 16620 41228
rect 16764 41210 16816 41216
rect 16868 41206 16896 41550
rect 17144 41274 17172 41618
rect 17500 41472 17552 41478
rect 17500 41414 17552 41420
rect 17132 41268 17184 41274
rect 17132 41210 17184 41216
rect 16856 41200 16908 41206
rect 16856 41142 16908 41148
rect 17144 40934 17172 41210
rect 17512 41002 17540 41414
rect 17604 41206 17632 41958
rect 17592 41200 17644 41206
rect 17592 41142 17644 41148
rect 17500 40996 17552 41002
rect 17500 40938 17552 40944
rect 17132 40928 17184 40934
rect 17132 40870 17184 40876
rect 17408 40928 17460 40934
rect 17408 40870 17460 40876
rect 17420 40730 17448 40870
rect 17408 40724 17460 40730
rect 17408 40666 17460 40672
rect 16856 40656 16908 40662
rect 16856 40598 16908 40604
rect 16868 40390 16896 40598
rect 17408 40452 17460 40458
rect 17408 40394 17460 40400
rect 16856 40384 16908 40390
rect 16856 40326 16908 40332
rect 17316 39976 17368 39982
rect 17316 39918 17368 39924
rect 16948 39840 17000 39846
rect 16948 39782 17000 39788
rect 16960 39574 16988 39782
rect 17328 39642 17356 39918
rect 17316 39636 17368 39642
rect 17316 39578 17368 39584
rect 16948 39568 17000 39574
rect 16948 39510 17000 39516
rect 17420 39438 17448 40394
rect 17696 40390 17724 42094
rect 17880 42022 17908 42298
rect 17972 42294 18000 42327
rect 17960 42288 18012 42294
rect 17960 42230 18012 42236
rect 18064 42226 18092 43318
rect 18156 43246 18184 44134
rect 18326 44024 18382 44033
rect 18326 43959 18328 43968
rect 18380 43959 18382 43968
rect 18328 43930 18380 43936
rect 18432 43654 18460 44474
rect 19708 44464 19760 44470
rect 19892 44464 19944 44470
rect 19760 44412 19892 44418
rect 19708 44406 19944 44412
rect 19524 44396 19576 44402
rect 19720 44390 19932 44406
rect 19524 44338 19576 44344
rect 18972 44192 19024 44198
rect 18972 44134 19024 44140
rect 18420 43648 18472 43654
rect 18420 43590 18472 43596
rect 18432 43314 18460 43590
rect 18420 43308 18472 43314
rect 18420 43250 18472 43256
rect 18144 43240 18196 43246
rect 18144 43182 18196 43188
rect 18052 42220 18104 42226
rect 18052 42162 18104 42168
rect 18328 42152 18380 42158
rect 17958 42120 18014 42129
rect 18328 42094 18380 42100
rect 17958 42055 17960 42064
rect 18012 42055 18014 42064
rect 17960 42026 18012 42032
rect 17868 42016 17920 42022
rect 17868 41958 17920 41964
rect 17972 41682 18000 42026
rect 17960 41676 18012 41682
rect 17960 41618 18012 41624
rect 18340 41614 18368 42094
rect 18432 41818 18460 43250
rect 18984 43178 19012 44134
rect 19340 43920 19392 43926
rect 19340 43862 19392 43868
rect 18972 43172 19024 43178
rect 18972 43114 19024 43120
rect 19352 42906 19380 43862
rect 19432 43852 19484 43858
rect 19432 43794 19484 43800
rect 19444 43654 19472 43794
rect 19432 43648 19484 43654
rect 19432 43590 19484 43596
rect 19536 43450 19564 44338
rect 19708 44328 19760 44334
rect 19708 44270 19760 44276
rect 19720 43654 19748 44270
rect 20720 44260 20772 44266
rect 20720 44202 20772 44208
rect 19800 44192 19852 44198
rect 19800 44134 19852 44140
rect 19708 43648 19760 43654
rect 19708 43590 19760 43596
rect 19524 43444 19576 43450
rect 19524 43386 19576 43392
rect 19340 42900 19392 42906
rect 19340 42842 19392 42848
rect 19352 42158 19380 42842
rect 19340 42152 19392 42158
rect 19340 42094 19392 42100
rect 19720 42022 19748 43590
rect 19812 42362 19840 44134
rect 20732 43994 20760 44202
rect 21180 44192 21232 44198
rect 21180 44134 21232 44140
rect 20720 43988 20772 43994
rect 20720 43930 20772 43936
rect 21088 43784 21140 43790
rect 21088 43726 21140 43732
rect 21100 43654 21128 43726
rect 20076 43648 20128 43654
rect 20076 43590 20128 43596
rect 20168 43648 20220 43654
rect 20168 43590 20220 43596
rect 21088 43648 21140 43654
rect 21088 43590 21140 43596
rect 20088 43382 20116 43590
rect 20076 43376 20128 43382
rect 20076 43318 20128 43324
rect 19984 43104 20036 43110
rect 19984 43046 20036 43052
rect 19996 42906 20024 43046
rect 19984 42900 20036 42906
rect 19984 42842 20036 42848
rect 20180 42566 20208 43590
rect 20536 43444 20588 43450
rect 20536 43386 20588 43392
rect 20442 43208 20498 43217
rect 20352 43172 20404 43178
rect 20442 43143 20498 43152
rect 20352 43114 20404 43120
rect 20364 42770 20392 43114
rect 20456 42906 20484 43143
rect 20548 42906 20576 43386
rect 21192 43178 21220 44134
rect 21180 43172 21232 43178
rect 21180 43114 21232 43120
rect 20444 42900 20496 42906
rect 20444 42842 20496 42848
rect 20536 42900 20588 42906
rect 20536 42842 20588 42848
rect 20352 42764 20404 42770
rect 20352 42706 20404 42712
rect 20168 42560 20220 42566
rect 20168 42502 20220 42508
rect 19800 42356 19852 42362
rect 19800 42298 19852 42304
rect 19708 42016 19760 42022
rect 19708 41958 19760 41964
rect 18420 41812 18472 41818
rect 18420 41754 18472 41760
rect 18788 41812 18840 41818
rect 18788 41754 18840 41760
rect 18328 41608 18380 41614
rect 18328 41550 18380 41556
rect 18420 41608 18472 41614
rect 18420 41550 18472 41556
rect 17960 41472 18012 41478
rect 17960 41414 18012 41420
rect 17868 41268 17920 41274
rect 17868 41210 17920 41216
rect 17776 40724 17828 40730
rect 17776 40666 17828 40672
rect 17684 40384 17736 40390
rect 17684 40326 17736 40332
rect 17408 39432 17460 39438
rect 17408 39374 17460 39380
rect 16764 38956 16816 38962
rect 16764 38898 16816 38904
rect 16488 37878 16540 37884
rect 16578 37904 16634 37913
rect 16578 37839 16634 37848
rect 16776 37330 16804 38898
rect 17592 38412 17644 38418
rect 17592 38354 17644 38360
rect 17684 38412 17736 38418
rect 17684 38354 17736 38360
rect 17604 38010 17632 38354
rect 17592 38004 17644 38010
rect 17592 37946 17644 37952
rect 17696 37466 17724 38354
rect 17788 37942 17816 40666
rect 17880 40390 17908 41210
rect 17868 40384 17920 40390
rect 17868 40326 17920 40332
rect 17880 38282 17908 40326
rect 17972 39846 18000 41414
rect 18328 40452 18380 40458
rect 18328 40394 18380 40400
rect 18340 40118 18368 40394
rect 18328 40112 18380 40118
rect 18328 40054 18380 40060
rect 17960 39840 18012 39846
rect 17960 39782 18012 39788
rect 18144 39840 18196 39846
rect 18144 39782 18196 39788
rect 18052 39500 18104 39506
rect 18052 39442 18104 39448
rect 18064 38758 18092 39442
rect 18052 38752 18104 38758
rect 18052 38694 18104 38700
rect 17868 38276 17920 38282
rect 17868 38218 17920 38224
rect 17776 37936 17828 37942
rect 17776 37878 17828 37884
rect 17868 37936 17920 37942
rect 17868 37878 17920 37884
rect 18064 37890 18092 38694
rect 18156 38010 18184 39782
rect 18432 39642 18460 41550
rect 18800 41138 18828 41754
rect 20180 41750 20208 42502
rect 20364 42072 20392 42706
rect 20456 42362 20484 42842
rect 20536 42696 20588 42702
rect 20536 42638 20588 42644
rect 20548 42566 20576 42638
rect 21284 42634 21312 44950
rect 27986 44840 28042 44849
rect 22836 44804 22888 44810
rect 27986 44775 28042 44784
rect 22836 44746 22888 44752
rect 21456 44736 21508 44742
rect 21456 44678 21508 44684
rect 22008 44736 22060 44742
rect 22008 44678 22060 44684
rect 21468 43722 21496 44678
rect 21640 44464 21692 44470
rect 21640 44406 21692 44412
rect 21548 43988 21600 43994
rect 21548 43930 21600 43936
rect 21456 43716 21508 43722
rect 21560 43704 21588 43930
rect 21652 43858 21680 44406
rect 22020 44402 22048 44678
rect 21916 44396 21968 44402
rect 21916 44338 21968 44344
rect 22008 44396 22060 44402
rect 22008 44338 22060 44344
rect 21732 44192 21784 44198
rect 21732 44134 21784 44140
rect 21744 43994 21772 44134
rect 21732 43988 21784 43994
rect 21732 43930 21784 43936
rect 21928 43926 21956 44338
rect 22560 44328 22612 44334
rect 22560 44270 22612 44276
rect 21916 43920 21968 43926
rect 21916 43862 21968 43868
rect 21640 43852 21692 43858
rect 21640 43794 21692 43800
rect 22284 43852 22336 43858
rect 22284 43794 22336 43800
rect 22100 43784 22152 43790
rect 22100 43726 22152 43732
rect 21824 43716 21876 43722
rect 21560 43676 21680 43704
rect 21456 43658 21508 43664
rect 21652 43178 21680 43676
rect 21824 43658 21876 43664
rect 21640 43172 21692 43178
rect 21640 43114 21692 43120
rect 21364 42696 21416 42702
rect 21362 42664 21364 42673
rect 21416 42664 21418 42673
rect 21272 42628 21324 42634
rect 21362 42599 21418 42608
rect 21272 42570 21324 42576
rect 20536 42560 20588 42566
rect 20536 42502 20588 42508
rect 20444 42356 20496 42362
rect 20444 42298 20496 42304
rect 20548 42226 20576 42502
rect 20536 42220 20588 42226
rect 20536 42162 20588 42168
rect 20444 42084 20496 42090
rect 20364 42044 20444 42072
rect 20444 42026 20496 42032
rect 21456 42084 21508 42090
rect 21456 42026 21508 42032
rect 20168 41744 20220 41750
rect 20168 41686 20220 41692
rect 19340 41676 19392 41682
rect 19340 41618 19392 41624
rect 19064 41540 19116 41546
rect 19064 41482 19116 41488
rect 18604 41132 18656 41138
rect 18604 41074 18656 41080
rect 18788 41132 18840 41138
rect 18788 41074 18840 41080
rect 18616 41018 18644 41074
rect 19076 41070 19104 41482
rect 19064 41064 19116 41070
rect 18616 40990 18828 41018
rect 19064 41006 19116 41012
rect 18696 40928 18748 40934
rect 18696 40870 18748 40876
rect 18512 40588 18564 40594
rect 18512 40530 18564 40536
rect 18524 40361 18552 40530
rect 18510 40352 18566 40361
rect 18510 40287 18566 40296
rect 18708 40186 18736 40870
rect 18800 40526 18828 40990
rect 19248 40588 19300 40594
rect 19248 40530 19300 40536
rect 18788 40520 18840 40526
rect 18788 40462 18840 40468
rect 18696 40180 18748 40186
rect 18696 40122 18748 40128
rect 18420 39636 18472 39642
rect 18420 39578 18472 39584
rect 18144 38004 18196 38010
rect 18144 37946 18196 37952
rect 17684 37460 17736 37466
rect 17684 37402 17736 37408
rect 16764 37324 16816 37330
rect 16764 37266 16816 37272
rect 12346 36680 12402 36689
rect 12346 36615 12402 36624
rect 16394 36680 16450 36689
rect 16394 36615 16450 36624
rect 11704 36576 11756 36582
rect 11704 36518 11756 36524
rect 8484 36508 8536 36514
rect 8484 36450 8536 36456
rect 8496 35737 8524 36450
rect 17880 36009 17908 37878
rect 18064 37862 18184 37890
rect 18156 37806 18184 37862
rect 18144 37800 18196 37806
rect 18050 37768 18106 37777
rect 18144 37742 18196 37748
rect 18050 37703 18106 37712
rect 17958 37632 18014 37641
rect 17958 37567 18014 37576
rect 17972 36553 18000 37567
rect 17958 36544 18014 36553
rect 17958 36479 18014 36488
rect 17866 36000 17922 36009
rect 17866 35935 17922 35944
rect 8206 35728 8262 35737
rect 8206 35663 8262 35672
rect 8482 35728 8538 35737
rect 8482 35663 8538 35672
rect 8220 35562 8248 35663
rect 18064 35562 18092 37703
rect 18156 37330 18184 37742
rect 18432 37466 18460 39578
rect 18512 39568 18564 39574
rect 18512 39510 18564 39516
rect 18524 37806 18552 39510
rect 18800 38350 18828 40462
rect 19064 39976 19116 39982
rect 19064 39918 19116 39924
rect 19076 39642 19104 39918
rect 19064 39636 19116 39642
rect 19064 39578 19116 39584
rect 19076 38962 19104 39578
rect 19064 38956 19116 38962
rect 19064 38898 19116 38904
rect 19260 38758 19288 40530
rect 19352 40390 19380 41618
rect 20180 41206 20208 41686
rect 20168 41200 20220 41206
rect 20168 41142 20220 41148
rect 19524 40996 19576 41002
rect 19524 40938 19576 40944
rect 19340 40384 19392 40390
rect 19340 40326 19392 40332
rect 19248 38752 19300 38758
rect 19248 38694 19300 38700
rect 19352 38554 19380 40326
rect 19536 38826 19564 40938
rect 20180 40934 20208 41142
rect 20168 40928 20220 40934
rect 20168 40870 20220 40876
rect 20456 39982 20484 42026
rect 21468 41478 21496 42026
rect 21272 41472 21324 41478
rect 21272 41414 21324 41420
rect 21456 41472 21508 41478
rect 21456 41414 21508 41420
rect 20720 40520 20772 40526
rect 20720 40462 20772 40468
rect 20810 40488 20866 40497
rect 20732 40186 20760 40462
rect 20810 40423 20866 40432
rect 20720 40180 20772 40186
rect 20720 40122 20772 40128
rect 20444 39976 20496 39982
rect 20444 39918 20496 39924
rect 20824 39522 20852 40423
rect 21284 39982 21312 41414
rect 21456 40520 21508 40526
rect 21456 40462 21508 40468
rect 21548 40520 21600 40526
rect 21548 40462 21600 40468
rect 21468 40390 21496 40462
rect 21456 40384 21508 40390
rect 21456 40326 21508 40332
rect 21468 40118 21496 40326
rect 21560 40186 21588 40462
rect 21652 40390 21680 43114
rect 21836 42090 21864 43658
rect 22008 43104 22060 43110
rect 22008 43046 22060 43052
rect 22020 42226 22048 43046
rect 22008 42220 22060 42226
rect 22008 42162 22060 42168
rect 21824 42084 21876 42090
rect 21824 42026 21876 42032
rect 21836 40662 21864 42026
rect 22020 41546 22048 42162
rect 22112 42158 22140 43726
rect 22192 42628 22244 42634
rect 22192 42570 22244 42576
rect 22100 42152 22152 42158
rect 22100 42094 22152 42100
rect 22098 41712 22154 41721
rect 22098 41647 22154 41656
rect 22112 41614 22140 41647
rect 22100 41608 22152 41614
rect 22100 41550 22152 41556
rect 22008 41540 22060 41546
rect 22008 41482 22060 41488
rect 22020 41414 22048 41482
rect 21928 41386 22048 41414
rect 21824 40656 21876 40662
rect 21824 40598 21876 40604
rect 21732 40520 21784 40526
rect 21732 40462 21784 40468
rect 21640 40384 21692 40390
rect 21640 40326 21692 40332
rect 21548 40180 21600 40186
rect 21548 40122 21600 40128
rect 21364 40112 21416 40118
rect 21364 40054 21416 40060
rect 21456 40112 21508 40118
rect 21456 40054 21508 40060
rect 21272 39976 21324 39982
rect 21272 39918 21324 39924
rect 21272 39840 21324 39846
rect 21272 39782 21324 39788
rect 21284 39642 21312 39782
rect 21376 39642 21404 40054
rect 21272 39636 21324 39642
rect 21272 39578 21324 39584
rect 21364 39636 21416 39642
rect 21364 39578 21416 39584
rect 20732 39494 20852 39522
rect 20536 39296 20588 39302
rect 20536 39238 20588 39244
rect 20168 39092 20220 39098
rect 20168 39034 20220 39040
rect 19524 38820 19576 38826
rect 19524 38762 19576 38768
rect 19616 38820 19668 38826
rect 19616 38762 19668 38768
rect 19340 38548 19392 38554
rect 19340 38490 19392 38496
rect 19248 38480 19300 38486
rect 19248 38422 19300 38428
rect 18788 38344 18840 38350
rect 18788 38286 18840 38292
rect 19260 38214 19288 38422
rect 19248 38208 19300 38214
rect 19248 38150 19300 38156
rect 19340 38208 19392 38214
rect 19340 38150 19392 38156
rect 18788 38004 18840 38010
rect 18788 37946 18840 37952
rect 18512 37800 18564 37806
rect 18512 37742 18564 37748
rect 18800 37670 18828 37946
rect 18788 37664 18840 37670
rect 18788 37606 18840 37612
rect 19064 37664 19116 37670
rect 19064 37606 19116 37612
rect 18420 37460 18472 37466
rect 18420 37402 18472 37408
rect 19076 37330 19104 37606
rect 18144 37324 18196 37330
rect 18144 37266 18196 37272
rect 19064 37324 19116 37330
rect 19064 37266 19116 37272
rect 19260 37262 19288 38150
rect 19352 38010 19380 38150
rect 19628 38010 19656 38762
rect 19340 38004 19392 38010
rect 19340 37946 19392 37952
rect 19616 38004 19668 38010
rect 19616 37946 19668 37952
rect 20180 37806 20208 39034
rect 20548 38554 20576 39238
rect 20536 38548 20588 38554
rect 20536 38490 20588 38496
rect 20732 38400 20760 39494
rect 20812 39432 20864 39438
rect 20812 39374 20864 39380
rect 20640 38372 20760 38400
rect 20640 38010 20668 38372
rect 20720 38276 20772 38282
rect 20720 38218 20772 38224
rect 20732 38010 20760 38218
rect 20628 38004 20680 38010
rect 20628 37946 20680 37952
rect 20720 38004 20772 38010
rect 20720 37946 20772 37952
rect 20168 37800 20220 37806
rect 20168 37742 20220 37748
rect 20824 37738 20852 39374
rect 21178 39264 21234 39273
rect 21178 39199 21234 39208
rect 21086 38992 21142 39001
rect 21086 38927 21142 38936
rect 20904 38208 20956 38214
rect 20904 38150 20956 38156
rect 20916 37738 20944 38150
rect 20996 38004 21048 38010
rect 20996 37946 21048 37952
rect 20812 37732 20864 37738
rect 20812 37674 20864 37680
rect 20904 37732 20956 37738
rect 20904 37674 20956 37680
rect 19340 37664 19392 37670
rect 19340 37606 19392 37612
rect 20260 37664 20312 37670
rect 20260 37606 20312 37612
rect 19248 37256 19300 37262
rect 19248 37198 19300 37204
rect 19352 36961 19380 37606
rect 20272 37466 20300 37606
rect 20260 37460 20312 37466
rect 20260 37402 20312 37408
rect 20720 37392 20772 37398
rect 20720 37334 20772 37340
rect 20628 37188 20680 37194
rect 20628 37130 20680 37136
rect 19338 36952 19394 36961
rect 19338 36887 19394 36896
rect 20076 35896 20128 35902
rect 20640 35873 20668 37130
rect 20732 36825 20760 37334
rect 20824 37262 20852 37674
rect 20812 37256 20864 37262
rect 20812 37198 20864 37204
rect 20718 36816 20774 36825
rect 20718 36751 20774 36760
rect 21008 36009 21036 37946
rect 21100 37233 21128 38927
rect 21086 37224 21142 37233
rect 21086 37159 21142 37168
rect 21192 37097 21220 39199
rect 21364 38752 21416 38758
rect 21364 38694 21416 38700
rect 21376 37738 21404 38694
rect 21468 38282 21496 40054
rect 21744 39914 21772 40462
rect 21824 40044 21876 40050
rect 21824 39986 21876 39992
rect 21732 39908 21784 39914
rect 21732 39850 21784 39856
rect 21744 39506 21772 39850
rect 21548 39500 21600 39506
rect 21548 39442 21600 39448
rect 21732 39500 21784 39506
rect 21732 39442 21784 39448
rect 21456 38276 21508 38282
rect 21456 38218 21508 38224
rect 21364 37732 21416 37738
rect 21364 37674 21416 37680
rect 21178 37088 21234 37097
rect 21178 37023 21234 37032
rect 21180 36848 21232 36854
rect 21180 36790 21232 36796
rect 20994 36000 21050 36009
rect 20994 35935 21050 35944
rect 20076 35838 20128 35844
rect 20626 35864 20682 35873
rect 20088 35737 20116 35838
rect 20626 35799 20682 35808
rect 21192 35737 21220 36790
rect 21560 36446 21588 39442
rect 21836 39438 21864 39986
rect 21824 39432 21876 39438
rect 21824 39374 21876 39380
rect 21732 39024 21784 39030
rect 21732 38966 21784 38972
rect 21744 38894 21772 38966
rect 21928 38962 21956 41386
rect 22008 40996 22060 41002
rect 22008 40938 22060 40944
rect 22020 40730 22048 40938
rect 22204 40934 22232 42570
rect 22296 42294 22324 43794
rect 22376 43784 22428 43790
rect 22376 43726 22428 43732
rect 22388 42566 22416 43726
rect 22468 43648 22520 43654
rect 22468 43590 22520 43596
rect 22376 42560 22428 42566
rect 22376 42502 22428 42508
rect 22284 42288 22336 42294
rect 22284 42230 22336 42236
rect 22284 42016 22336 42022
rect 22284 41958 22336 41964
rect 22192 40928 22244 40934
rect 22192 40870 22244 40876
rect 22008 40724 22060 40730
rect 22008 40666 22060 40672
rect 22204 40458 22232 40870
rect 22192 40452 22244 40458
rect 22192 40394 22244 40400
rect 22008 40384 22060 40390
rect 22008 40326 22060 40332
rect 21916 38956 21968 38962
rect 21916 38898 21968 38904
rect 21732 38888 21784 38894
rect 21732 38830 21784 38836
rect 21640 38548 21692 38554
rect 21744 38536 21772 38830
rect 21692 38508 21772 38536
rect 21640 38490 21692 38496
rect 21928 38486 21956 38898
rect 22020 38758 22048 40326
rect 22204 38962 22232 40394
rect 22296 40050 22324 41958
rect 22388 41721 22416 42502
rect 22480 41818 22508 43590
rect 22572 43450 22600 44270
rect 22744 43784 22796 43790
rect 22744 43726 22796 43732
rect 22560 43444 22612 43450
rect 22560 43386 22612 43392
rect 22572 42770 22600 43386
rect 22652 42832 22704 42838
rect 22652 42774 22704 42780
rect 22560 42764 22612 42770
rect 22560 42706 22612 42712
rect 22560 42560 22612 42566
rect 22560 42502 22612 42508
rect 22572 42226 22600 42502
rect 22560 42220 22612 42226
rect 22560 42162 22612 42168
rect 22468 41812 22520 41818
rect 22468 41754 22520 41760
rect 22374 41712 22430 41721
rect 22374 41647 22430 41656
rect 22376 41608 22428 41614
rect 22376 41550 22428 41556
rect 22560 41608 22612 41614
rect 22560 41550 22612 41556
rect 22388 41478 22416 41550
rect 22376 41472 22428 41478
rect 22376 41414 22428 41420
rect 22284 40044 22336 40050
rect 22284 39986 22336 39992
rect 22572 39420 22600 41550
rect 22664 40905 22692 42774
rect 22756 42022 22784 43726
rect 22848 43110 22876 44746
rect 23296 44736 23348 44742
rect 23296 44678 23348 44684
rect 26424 44736 26476 44742
rect 26424 44678 26476 44684
rect 27342 44704 27398 44713
rect 23020 44464 23072 44470
rect 23020 44406 23072 44412
rect 23032 43926 23060 44406
rect 23020 43920 23072 43926
rect 23020 43862 23072 43868
rect 23308 43382 23336 44678
rect 24596 44526 25084 44554
rect 26436 44538 26464 44678
rect 27342 44639 27398 44648
rect 23480 44192 23532 44198
rect 23480 44134 23532 44140
rect 23664 44192 23716 44198
rect 23664 44134 23716 44140
rect 24216 44192 24268 44198
rect 24216 44134 24268 44140
rect 23388 43784 23440 43790
rect 23388 43726 23440 43732
rect 23400 43450 23428 43726
rect 23388 43444 23440 43450
rect 23388 43386 23440 43392
rect 23296 43376 23348 43382
rect 23296 43318 23348 43324
rect 22836 43104 22888 43110
rect 22836 43046 22888 43052
rect 23020 43104 23072 43110
rect 23020 43046 23072 43052
rect 22848 42838 22876 43046
rect 22836 42832 22888 42838
rect 22836 42774 22888 42780
rect 22848 42566 22876 42774
rect 22836 42560 22888 42566
rect 22836 42502 22888 42508
rect 22744 42016 22796 42022
rect 22744 41958 22796 41964
rect 22848 41018 22876 42502
rect 23032 42158 23060 43046
rect 23308 42888 23336 43318
rect 23492 43246 23520 44134
rect 23676 43926 23704 44134
rect 23664 43920 23716 43926
rect 23664 43862 23716 43868
rect 23480 43240 23532 43246
rect 23480 43182 23532 43188
rect 23664 43240 23716 43246
rect 23664 43182 23716 43188
rect 23492 42906 23520 43182
rect 23216 42860 23336 42888
rect 23480 42900 23532 42906
rect 23020 42152 23072 42158
rect 23020 42094 23072 42100
rect 23110 41712 23166 41721
rect 23110 41647 23166 41656
rect 22848 40990 22968 41018
rect 22650 40896 22706 40905
rect 22650 40831 22706 40840
rect 22652 40588 22704 40594
rect 22652 40530 22704 40536
rect 22664 40050 22692 40530
rect 22744 40384 22796 40390
rect 22744 40326 22796 40332
rect 22652 40044 22704 40050
rect 22652 39986 22704 39992
rect 22756 39642 22784 40326
rect 22940 40118 22968 40990
rect 23020 40996 23072 41002
rect 23020 40938 23072 40944
rect 23032 40730 23060 40938
rect 23020 40724 23072 40730
rect 23020 40666 23072 40672
rect 23032 40458 23060 40666
rect 23020 40452 23072 40458
rect 23020 40394 23072 40400
rect 22928 40112 22980 40118
rect 22928 40054 22980 40060
rect 22744 39636 22796 39642
rect 22744 39578 22796 39584
rect 22652 39432 22704 39438
rect 22572 39392 22652 39420
rect 22652 39374 22704 39380
rect 22468 39364 22520 39370
rect 22468 39306 22520 39312
rect 22192 38956 22244 38962
rect 22192 38898 22244 38904
rect 22192 38820 22244 38826
rect 22192 38762 22244 38768
rect 22008 38752 22060 38758
rect 22008 38694 22060 38700
rect 22204 38554 22232 38762
rect 22100 38548 22152 38554
rect 22100 38490 22152 38496
rect 22192 38548 22244 38554
rect 22192 38490 22244 38496
rect 21916 38480 21968 38486
rect 21916 38422 21968 38428
rect 22112 38434 22140 38490
rect 22480 38434 22508 39306
rect 22112 38418 22508 38434
rect 22112 38412 22520 38418
rect 22112 38406 22468 38412
rect 22468 38354 22520 38360
rect 21732 38344 21784 38350
rect 21732 38286 21784 38292
rect 21744 37670 21772 38286
rect 21732 37664 21784 37670
rect 21732 37606 21784 37612
rect 21744 37466 21772 37606
rect 21732 37460 21784 37466
rect 21732 37402 21784 37408
rect 22008 36780 22060 36786
rect 22008 36722 22060 36728
rect 21548 36440 21600 36446
rect 21548 36382 21600 36388
rect 22020 35737 22048 36722
rect 23124 35902 23152 41647
rect 23216 40662 23244 42860
rect 23480 42842 23532 42848
rect 23296 42016 23348 42022
rect 23296 41958 23348 41964
rect 23308 41750 23336 41958
rect 23296 41744 23348 41750
rect 23296 41686 23348 41692
rect 23296 41472 23348 41478
rect 23296 41414 23348 41420
rect 23308 41206 23336 41414
rect 23296 41200 23348 41206
rect 23296 41142 23348 41148
rect 23204 40656 23256 40662
rect 23204 40598 23256 40604
rect 23308 40050 23336 41142
rect 23296 40044 23348 40050
rect 23296 39986 23348 39992
rect 23492 39982 23520 42842
rect 23676 41818 23704 43182
rect 24228 43178 24256 44134
rect 24216 43172 24268 43178
rect 24216 43114 24268 43120
rect 24596 42684 24624 44526
rect 25056 44402 25084 44526
rect 26332 44532 26384 44538
rect 26332 44474 26384 44480
rect 26424 44532 26476 44538
rect 26424 44474 26476 44480
rect 25686 44432 25742 44441
rect 24768 44396 24820 44402
rect 25044 44396 25096 44402
rect 24820 44356 24992 44384
rect 24768 44338 24820 44344
rect 24676 44192 24728 44198
rect 24676 44134 24728 44140
rect 24768 44192 24820 44198
rect 24768 44134 24820 44140
rect 24688 43994 24716 44134
rect 24676 43988 24728 43994
rect 24676 43930 24728 43936
rect 24676 42696 24728 42702
rect 24214 42664 24270 42673
rect 24214 42599 24270 42608
rect 24596 42656 24676 42684
rect 24228 42566 24256 42599
rect 24216 42560 24268 42566
rect 24216 42502 24268 42508
rect 24032 42220 24084 42226
rect 24032 42162 24084 42168
rect 23756 42152 23808 42158
rect 23756 42094 23808 42100
rect 23664 41812 23716 41818
rect 23664 41754 23716 41760
rect 23768 41206 23796 42094
rect 24044 41614 24072 42162
rect 24032 41608 24084 41614
rect 24032 41550 24084 41556
rect 24596 41414 24624 42656
rect 24676 42638 24728 42644
rect 24780 42362 24808 44134
rect 24964 43994 24992 44356
rect 25686 44367 25688 44376
rect 25044 44338 25096 44344
rect 25740 44367 25742 44376
rect 25688 44338 25740 44344
rect 25228 44260 25280 44266
rect 25228 44202 25280 44208
rect 25504 44260 25556 44266
rect 25504 44202 25556 44208
rect 24952 43988 25004 43994
rect 24952 43930 25004 43936
rect 24860 43920 24912 43926
rect 24860 43862 24912 43868
rect 24872 43178 24900 43862
rect 25240 43382 25268 44202
rect 25228 43376 25280 43382
rect 25228 43318 25280 43324
rect 24860 43172 24912 43178
rect 24860 43114 24912 43120
rect 24872 42838 24900 43114
rect 25412 43104 25464 43110
rect 24950 43072 25006 43081
rect 25516 43081 25544 44202
rect 25688 44192 25740 44198
rect 25688 44134 25740 44140
rect 25412 43046 25464 43052
rect 25502 43072 25558 43081
rect 24950 43007 25006 43016
rect 24964 42906 24992 43007
rect 24952 42900 25004 42906
rect 24952 42842 25004 42848
rect 24860 42832 24912 42838
rect 24860 42774 24912 42780
rect 24768 42356 24820 42362
rect 24768 42298 24820 42304
rect 24872 41682 24900 42774
rect 25044 42764 25096 42770
rect 25044 42706 25096 42712
rect 24952 42628 25004 42634
rect 24952 42570 25004 42576
rect 24964 42362 24992 42570
rect 24952 42356 25004 42362
rect 24952 42298 25004 42304
rect 25056 42158 25084 42706
rect 25136 42696 25188 42702
rect 25136 42638 25188 42644
rect 25228 42696 25280 42702
rect 25228 42638 25280 42644
rect 25318 42664 25374 42673
rect 25044 42152 25096 42158
rect 25044 42094 25096 42100
rect 25148 41818 25176 42638
rect 25240 42294 25268 42638
rect 25318 42599 25374 42608
rect 25228 42288 25280 42294
rect 25228 42230 25280 42236
rect 25226 41984 25282 41993
rect 25226 41919 25282 41928
rect 25136 41812 25188 41818
rect 25136 41754 25188 41760
rect 24860 41676 24912 41682
rect 24860 41618 24912 41624
rect 24674 41576 24730 41585
rect 24674 41511 24730 41520
rect 24504 41386 24624 41414
rect 23756 41200 23808 41206
rect 23756 41142 23808 41148
rect 24504 41138 24532 41386
rect 24492 41132 24544 41138
rect 24492 41074 24544 41080
rect 23756 40928 23808 40934
rect 23756 40870 23808 40876
rect 23768 40662 23796 40870
rect 23756 40656 23808 40662
rect 23756 40598 23808 40604
rect 23480 39976 23532 39982
rect 23480 39918 23532 39924
rect 24032 39976 24084 39982
rect 24032 39918 24084 39924
rect 23848 39840 23900 39846
rect 23848 39782 23900 39788
rect 23388 38956 23440 38962
rect 23388 38898 23440 38904
rect 23400 37806 23428 38898
rect 23860 38554 23888 39782
rect 24044 39642 24072 39918
rect 24032 39636 24084 39642
rect 24032 39578 24084 39584
rect 24044 39250 24072 39578
rect 24308 39432 24360 39438
rect 24308 39374 24360 39380
rect 23952 39222 24072 39250
rect 24124 39296 24176 39302
rect 24124 39238 24176 39244
rect 23952 39098 23980 39222
rect 23940 39092 23992 39098
rect 23940 39034 23992 39040
rect 24136 38962 24164 39238
rect 24320 39098 24348 39374
rect 24308 39092 24360 39098
rect 24308 39034 24360 39040
rect 24124 38956 24176 38962
rect 24124 38898 24176 38904
rect 24216 38956 24268 38962
rect 24216 38898 24268 38904
rect 23848 38548 23900 38554
rect 23848 38490 23900 38496
rect 23572 38344 23624 38350
rect 23572 38286 23624 38292
rect 24032 38344 24084 38350
rect 24228 38332 24256 38898
rect 24084 38304 24256 38332
rect 24032 38286 24084 38292
rect 23584 38010 23612 38286
rect 23572 38004 23624 38010
rect 23572 37946 23624 37952
rect 23388 37800 23440 37806
rect 23388 37742 23440 37748
rect 24216 37664 24268 37670
rect 24320 37652 24348 39034
rect 24504 38962 24532 41074
rect 24688 41002 24716 41511
rect 24872 41478 24900 41618
rect 24860 41472 24912 41478
rect 24860 41414 24912 41420
rect 24676 40996 24728 41002
rect 24676 40938 24728 40944
rect 24768 40996 24820 41002
rect 24768 40938 24820 40944
rect 24688 39574 24716 40938
rect 24780 40526 24808 40938
rect 24768 40520 24820 40526
rect 24872 40508 24900 41414
rect 25136 40928 25188 40934
rect 25136 40870 25188 40876
rect 24952 40520 25004 40526
rect 24872 40480 24952 40508
rect 24768 40462 24820 40468
rect 24952 40462 25004 40468
rect 24964 39914 24992 40462
rect 25044 40452 25096 40458
rect 25044 40394 25096 40400
rect 25056 40089 25084 40394
rect 25042 40080 25098 40089
rect 25042 40015 25098 40024
rect 24860 39908 24912 39914
rect 24860 39850 24912 39856
rect 24952 39908 25004 39914
rect 24952 39850 25004 39856
rect 24872 39574 24900 39850
rect 24676 39568 24728 39574
rect 24676 39510 24728 39516
rect 24860 39568 24912 39574
rect 24860 39510 24912 39516
rect 24492 38956 24544 38962
rect 24492 38898 24544 38904
rect 24964 38758 24992 39850
rect 25148 39642 25176 40870
rect 25136 39636 25188 39642
rect 25136 39578 25188 39584
rect 25042 39536 25098 39545
rect 25042 39471 25098 39480
rect 25056 39273 25084 39471
rect 25042 39264 25098 39273
rect 25042 39199 25098 39208
rect 24952 38752 25004 38758
rect 24952 38694 25004 38700
rect 24582 38584 24638 38593
rect 24582 38519 24584 38528
rect 24636 38519 24638 38528
rect 24584 38490 24636 38496
rect 25044 38480 25096 38486
rect 25044 38422 25096 38428
rect 25056 37738 25084 38422
rect 24952 37732 25004 37738
rect 24952 37674 25004 37680
rect 25044 37732 25096 37738
rect 25044 37674 25096 37680
rect 24268 37624 24348 37652
rect 24860 37664 24912 37670
rect 24216 37606 24268 37612
rect 24860 37606 24912 37612
rect 23204 37324 23256 37330
rect 23204 37266 23256 37272
rect 23216 36825 23244 37266
rect 23478 37224 23534 37233
rect 23478 37159 23534 37168
rect 23492 36922 23520 37159
rect 23480 36916 23532 36922
rect 23480 36858 23532 36864
rect 23202 36816 23258 36825
rect 23202 36751 23258 36760
rect 24872 36650 24900 37606
rect 24964 37466 24992 37674
rect 24952 37460 25004 37466
rect 24952 37402 25004 37408
rect 25056 37330 25084 37674
rect 25044 37324 25096 37330
rect 25044 37266 25096 37272
rect 25240 37194 25268 41919
rect 25332 41414 25360 42599
rect 25424 42022 25452 43046
rect 25502 43007 25558 43016
rect 25700 42702 25728 44134
rect 26240 43852 26292 43858
rect 26240 43794 26292 43800
rect 25872 43648 25924 43654
rect 26056 43648 26108 43654
rect 25872 43590 25924 43596
rect 25962 43616 26018 43625
rect 25780 43444 25832 43450
rect 25780 43386 25832 43392
rect 25792 42906 25820 43386
rect 25884 43110 25912 43590
rect 26056 43590 26108 43596
rect 25962 43551 26018 43560
rect 25872 43104 25924 43110
rect 25872 43046 25924 43052
rect 25976 42906 26004 43551
rect 26068 43246 26096 43590
rect 26252 43314 26280 43794
rect 26240 43308 26292 43314
rect 26240 43250 26292 43256
rect 26056 43240 26108 43246
rect 26056 43182 26108 43188
rect 25780 42900 25832 42906
rect 25780 42842 25832 42848
rect 25964 42900 26016 42906
rect 25964 42842 26016 42848
rect 25688 42696 25740 42702
rect 25688 42638 25740 42644
rect 25412 42016 25464 42022
rect 25412 41958 25464 41964
rect 25502 41848 25558 41857
rect 25502 41783 25558 41792
rect 25332 41386 25452 41414
rect 25320 40384 25372 40390
rect 25320 40326 25372 40332
rect 25332 40186 25360 40326
rect 25320 40180 25372 40186
rect 25320 40122 25372 40128
rect 25228 37188 25280 37194
rect 25228 37130 25280 37136
rect 24860 36644 24912 36650
rect 24860 36586 24912 36592
rect 25424 36145 25452 41386
rect 25410 36136 25466 36145
rect 23204 36100 23256 36106
rect 25410 36071 25466 36080
rect 23204 36042 23256 36048
rect 23112 35896 23164 35902
rect 23216 35873 23244 36042
rect 24676 36032 24728 36038
rect 24674 36000 24676 36009
rect 24728 36000 24730 36009
rect 24674 35935 24730 35944
rect 23572 35896 23624 35902
rect 23112 35838 23164 35844
rect 23202 35864 23258 35873
rect 25516 35873 25544 41783
rect 25700 41614 25728 42638
rect 25976 42362 26004 42842
rect 26068 42770 26096 43182
rect 26240 43104 26292 43110
rect 26240 43046 26292 43052
rect 26146 42936 26202 42945
rect 26252 42906 26280 43046
rect 26344 42906 26372 44474
rect 27356 44402 27384 44639
rect 27344 44396 27396 44402
rect 27344 44338 27396 44344
rect 28000 44334 28028 44775
rect 29092 44736 29144 44742
rect 28722 44704 28778 44713
rect 29092 44678 29144 44684
rect 32404 44736 32456 44742
rect 32404 44678 32456 44684
rect 28722 44639 28778 44648
rect 28736 44402 28764 44639
rect 28080 44396 28132 44402
rect 28080 44338 28132 44344
rect 28724 44396 28776 44402
rect 28724 44338 28776 44344
rect 27988 44328 28040 44334
rect 27988 44270 28040 44276
rect 26884 44260 26936 44266
rect 26884 44202 26936 44208
rect 26516 44192 26568 44198
rect 26516 44134 26568 44140
rect 26424 43376 26476 43382
rect 26424 43318 26476 43324
rect 26146 42871 26202 42880
rect 26240 42900 26292 42906
rect 26056 42764 26108 42770
rect 26056 42706 26108 42712
rect 25964 42356 26016 42362
rect 25964 42298 26016 42304
rect 25780 42016 25832 42022
rect 25780 41958 25832 41964
rect 25792 41721 25820 41958
rect 25778 41712 25834 41721
rect 25778 41647 25834 41656
rect 26054 41712 26110 41721
rect 26054 41647 26110 41656
rect 25688 41608 25740 41614
rect 25688 41550 25740 41556
rect 25964 41608 26016 41614
rect 25964 41550 26016 41556
rect 25870 41304 25926 41313
rect 25870 41239 25926 41248
rect 25596 39432 25648 39438
rect 25596 39374 25648 39380
rect 25608 39030 25636 39374
rect 25596 39024 25648 39030
rect 25596 38966 25648 38972
rect 25688 38752 25740 38758
rect 25688 38694 25740 38700
rect 25700 38350 25728 38694
rect 25688 38344 25740 38350
rect 25884 38298 25912 41239
rect 25976 41041 26004 41550
rect 26068 41449 26096 41647
rect 26054 41440 26110 41449
rect 26054 41375 26110 41384
rect 26160 41041 26188 42871
rect 26240 42842 26292 42848
rect 26332 42900 26384 42906
rect 26332 42842 26384 42848
rect 26436 41682 26464 43318
rect 26528 42770 26556 44134
rect 26896 43858 26924 44202
rect 27896 44192 27948 44198
rect 27896 44134 27948 44140
rect 27908 43926 27936 44134
rect 27896 43920 27948 43926
rect 27896 43862 27948 43868
rect 26884 43852 26936 43858
rect 26884 43794 26936 43800
rect 26792 43784 26844 43790
rect 26792 43726 26844 43732
rect 27252 43784 27304 43790
rect 27252 43726 27304 43732
rect 26608 43716 26660 43722
rect 26608 43658 26660 43664
rect 26516 42764 26568 42770
rect 26516 42706 26568 42712
rect 26516 42628 26568 42634
rect 26516 42570 26568 42576
rect 26240 41676 26292 41682
rect 26240 41618 26292 41624
rect 26424 41676 26476 41682
rect 26424 41618 26476 41624
rect 25962 41032 26018 41041
rect 25962 40967 26018 40976
rect 26146 41032 26202 41041
rect 26146 40967 26202 40976
rect 26252 40934 26280 41618
rect 26528 41414 26556 42570
rect 26620 42226 26648 43658
rect 26700 42560 26752 42566
rect 26700 42502 26752 42508
rect 26608 42220 26660 42226
rect 26608 42162 26660 42168
rect 26436 41386 26556 41414
rect 26240 40928 26292 40934
rect 26240 40870 26292 40876
rect 26252 40730 26280 40870
rect 26240 40724 26292 40730
rect 26240 40666 26292 40672
rect 26056 40520 26108 40526
rect 26056 40462 26108 40468
rect 26068 39370 26096 40462
rect 26252 39982 26280 40666
rect 26240 39976 26292 39982
rect 26240 39918 26292 39924
rect 26056 39364 26108 39370
rect 26056 39306 26108 39312
rect 25964 39296 26016 39302
rect 25964 39238 26016 39244
rect 25688 38286 25740 38292
rect 25792 38270 25912 38298
rect 25792 37505 25820 38270
rect 25872 38208 25924 38214
rect 25872 38150 25924 38156
rect 25778 37496 25834 37505
rect 25884 37466 25912 38150
rect 25976 37466 26004 39238
rect 26068 39098 26096 39306
rect 26056 39092 26108 39098
rect 26056 39034 26108 39040
rect 26148 38752 26200 38758
rect 26148 38694 26200 38700
rect 26160 37466 26188 38694
rect 26252 38554 26280 39918
rect 26332 39840 26384 39846
rect 26332 39782 26384 39788
rect 26344 39642 26372 39782
rect 26332 39636 26384 39642
rect 26332 39578 26384 39584
rect 26436 39522 26464 41386
rect 26620 41138 26648 42162
rect 26712 41750 26740 42502
rect 26700 41744 26752 41750
rect 26700 41686 26752 41692
rect 26804 41206 26832 43726
rect 26884 42560 26936 42566
rect 26884 42502 26936 42508
rect 26896 42090 26924 42502
rect 26884 42084 26936 42090
rect 26884 42026 26936 42032
rect 26792 41200 26844 41206
rect 26792 41142 26844 41148
rect 26608 41132 26660 41138
rect 26528 41092 26608 41120
rect 26528 40730 26556 41092
rect 26608 41074 26660 41080
rect 26516 40724 26568 40730
rect 26516 40666 26568 40672
rect 26528 40050 26556 40666
rect 27264 40662 27292 43726
rect 28092 43382 28120 44338
rect 28816 44192 28868 44198
rect 28816 44134 28868 44140
rect 28828 43450 28856 44134
rect 29104 43926 29132 44678
rect 32416 44538 32444 44678
rect 32404 44532 32456 44538
rect 32404 44474 32456 44480
rect 32956 44532 33008 44538
rect 32956 44474 33008 44480
rect 31024 44328 31076 44334
rect 31024 44270 31076 44276
rect 29092 43920 29144 43926
rect 29092 43862 29144 43868
rect 28816 43444 28868 43450
rect 28816 43386 28868 43392
rect 28908 43444 28960 43450
rect 28908 43386 28960 43392
rect 27436 43376 27488 43382
rect 27436 43318 27488 43324
rect 28080 43376 28132 43382
rect 28080 43318 28132 43324
rect 27448 43110 27476 43318
rect 27528 43172 27580 43178
rect 27528 43114 27580 43120
rect 27344 43104 27396 43110
rect 27344 43046 27396 43052
rect 27436 43104 27488 43110
rect 27436 43046 27488 43052
rect 27356 42906 27384 43046
rect 27344 42900 27396 42906
rect 27344 42842 27396 42848
rect 27540 42770 27568 43114
rect 27988 42900 28040 42906
rect 27988 42842 28040 42848
rect 27528 42764 27580 42770
rect 27528 42706 27580 42712
rect 27436 42220 27488 42226
rect 27436 42162 27488 42168
rect 27448 41818 27476 42162
rect 27436 41812 27488 41818
rect 27436 41754 27488 41760
rect 27620 41812 27672 41818
rect 27620 41754 27672 41760
rect 27632 41562 27660 41754
rect 27356 41534 27660 41562
rect 27356 41478 27384 41534
rect 27344 41472 27396 41478
rect 27344 41414 27396 41420
rect 28000 41274 28028 42842
rect 28092 42702 28120 43318
rect 28540 43308 28592 43314
rect 28540 43250 28592 43256
rect 28356 43240 28408 43246
rect 28356 43182 28408 43188
rect 28080 42696 28132 42702
rect 28080 42638 28132 42644
rect 28368 42684 28396 43182
rect 28552 42770 28580 43250
rect 28920 43178 28948 43386
rect 28908 43172 28960 43178
rect 28908 43114 28960 43120
rect 28540 42764 28592 42770
rect 28540 42706 28592 42712
rect 28448 42696 28500 42702
rect 28368 42656 28448 42684
rect 28092 42294 28120 42638
rect 28368 42362 28396 42656
rect 28448 42638 28500 42644
rect 28356 42356 28408 42362
rect 28356 42298 28408 42304
rect 28080 42288 28132 42294
rect 28080 42230 28132 42236
rect 28816 42288 28868 42294
rect 28816 42230 28868 42236
rect 28448 42152 28500 42158
rect 28448 42094 28500 42100
rect 28264 42016 28316 42022
rect 28264 41958 28316 41964
rect 28276 41750 28304 41958
rect 28264 41744 28316 41750
rect 28264 41686 28316 41692
rect 28264 41540 28316 41546
rect 28264 41482 28316 41488
rect 28356 41540 28408 41546
rect 28356 41482 28408 41488
rect 27988 41268 28040 41274
rect 27988 41210 28040 41216
rect 28276 40730 28304 41482
rect 28368 41070 28396 41482
rect 28356 41064 28408 41070
rect 28356 41006 28408 41012
rect 27436 40724 27488 40730
rect 27436 40666 27488 40672
rect 28264 40724 28316 40730
rect 28264 40666 28316 40672
rect 27252 40656 27304 40662
rect 27252 40598 27304 40604
rect 27068 40520 27120 40526
rect 27068 40462 27120 40468
rect 26608 40384 26660 40390
rect 26608 40326 26660 40332
rect 26516 40044 26568 40050
rect 26516 39986 26568 39992
rect 26344 39494 26464 39522
rect 26240 38548 26292 38554
rect 26240 38490 26292 38496
rect 26252 37874 26280 38490
rect 26344 38010 26372 39494
rect 26424 39432 26476 39438
rect 26424 39374 26476 39380
rect 26332 38004 26384 38010
rect 26332 37946 26384 37952
rect 26240 37868 26292 37874
rect 26240 37810 26292 37816
rect 26332 37732 26384 37738
rect 26332 37674 26384 37680
rect 25778 37431 25834 37440
rect 25872 37460 25924 37466
rect 25872 37402 25924 37408
rect 25964 37460 26016 37466
rect 25964 37402 26016 37408
rect 26148 37460 26200 37466
rect 26148 37402 26200 37408
rect 26344 37330 26372 37674
rect 26436 37670 26464 39374
rect 26516 39296 26568 39302
rect 26516 39238 26568 39244
rect 26528 38894 26556 39238
rect 26516 38888 26568 38894
rect 26516 38830 26568 38836
rect 26620 38729 26648 40326
rect 27080 39846 27108 40462
rect 27448 40186 27476 40666
rect 27528 40452 27580 40458
rect 27528 40394 27580 40400
rect 27540 40186 27568 40394
rect 27436 40180 27488 40186
rect 27436 40122 27488 40128
rect 27528 40180 27580 40186
rect 27528 40122 27580 40128
rect 27160 40044 27212 40050
rect 27160 39986 27212 39992
rect 27068 39840 27120 39846
rect 27068 39782 27120 39788
rect 26700 39024 26752 39030
rect 26700 38966 26752 38972
rect 26712 38894 26740 38966
rect 26700 38888 26752 38894
rect 26700 38830 26752 38836
rect 26792 38752 26844 38758
rect 26606 38720 26662 38729
rect 26792 38694 26844 38700
rect 26606 38655 26662 38664
rect 26698 38176 26754 38185
rect 26698 38111 26754 38120
rect 26516 38004 26568 38010
rect 26516 37946 26568 37952
rect 26424 37664 26476 37670
rect 26424 37606 26476 37612
rect 26436 37330 26464 37606
rect 26332 37324 26384 37330
rect 26332 37266 26384 37272
rect 26424 37324 26476 37330
rect 26424 37266 26476 37272
rect 26528 37262 26556 37946
rect 26712 37777 26740 38111
rect 26804 37874 26832 38694
rect 26976 38480 27028 38486
rect 26976 38422 27028 38428
rect 26792 37868 26844 37874
rect 26792 37810 26844 37816
rect 26698 37768 26754 37777
rect 26698 37703 26754 37712
rect 26516 37256 26568 37262
rect 26516 37198 26568 37204
rect 26988 37126 27016 38422
rect 27068 38344 27120 38350
rect 27172 38332 27200 39986
rect 27436 39840 27488 39846
rect 27436 39782 27488 39788
rect 28356 39840 28408 39846
rect 28356 39782 28408 39788
rect 27252 39296 27304 39302
rect 27252 39238 27304 39244
rect 27120 38304 27200 38332
rect 27068 38286 27120 38292
rect 27172 37874 27200 38304
rect 27160 37868 27212 37874
rect 27160 37810 27212 37816
rect 26976 37120 27028 37126
rect 26976 37062 27028 37068
rect 27264 36417 27292 39238
rect 27448 38593 27476 39782
rect 27618 39672 27674 39681
rect 28368 39642 28396 39782
rect 27618 39607 27674 39616
rect 28356 39636 28408 39642
rect 27632 39574 27660 39607
rect 28356 39578 28408 39584
rect 27620 39568 27672 39574
rect 27620 39510 27672 39516
rect 27620 39364 27672 39370
rect 27620 39306 27672 39312
rect 27896 39364 27948 39370
rect 27896 39306 27948 39312
rect 27632 39250 27660 39306
rect 27540 39222 27660 39250
rect 27434 38584 27490 38593
rect 27434 38519 27490 38528
rect 27448 37466 27476 38519
rect 27540 38214 27568 39222
rect 27632 38814 27844 38842
rect 27632 38486 27660 38814
rect 27816 38758 27844 38814
rect 27712 38752 27764 38758
rect 27712 38694 27764 38700
rect 27804 38752 27856 38758
rect 27804 38694 27856 38700
rect 27620 38480 27672 38486
rect 27620 38422 27672 38428
rect 27528 38208 27580 38214
rect 27528 38150 27580 38156
rect 27526 37632 27582 37641
rect 27526 37567 27582 37576
rect 27436 37460 27488 37466
rect 27436 37402 27488 37408
rect 27540 37194 27568 37567
rect 27724 37466 27752 38694
rect 27804 38004 27856 38010
rect 27804 37946 27856 37952
rect 27816 37913 27844 37946
rect 27802 37904 27858 37913
rect 27802 37839 27858 37848
rect 27712 37460 27764 37466
rect 27712 37402 27764 37408
rect 27528 37188 27580 37194
rect 27528 37130 27580 37136
rect 27908 36768 27936 39306
rect 27988 39092 28040 39098
rect 27988 39034 28040 39040
rect 28000 39001 28028 39034
rect 27986 38992 28042 39001
rect 27986 38927 28042 38936
rect 28264 38752 28316 38758
rect 28264 38694 28316 38700
rect 28276 37942 28304 38694
rect 28460 38418 28488 42094
rect 28724 41744 28776 41750
rect 28644 41704 28724 41732
rect 28538 38448 28594 38457
rect 28448 38412 28500 38418
rect 28538 38383 28594 38392
rect 28448 38354 28500 38360
rect 28356 38276 28408 38282
rect 28356 38218 28408 38224
rect 28368 38185 28396 38218
rect 28354 38176 28410 38185
rect 28354 38111 28410 38120
rect 28264 37936 28316 37942
rect 28264 37878 28316 37884
rect 28276 37806 28304 37878
rect 28264 37800 28316 37806
rect 28078 37768 28134 37777
rect 28264 37742 28316 37748
rect 28354 37768 28410 37777
rect 28078 37703 28080 37712
rect 28132 37703 28134 37712
rect 28354 37703 28410 37712
rect 28080 37674 28132 37680
rect 28368 37505 28396 37703
rect 28460 37670 28488 38354
rect 28552 38185 28580 38383
rect 28538 38176 28594 38185
rect 28538 38111 28594 38120
rect 28448 37664 28500 37670
rect 28448 37606 28500 37612
rect 28354 37496 28410 37505
rect 28354 37431 28410 37440
rect 28538 37496 28594 37505
rect 28538 37431 28594 37440
rect 27540 36740 27936 36768
rect 27540 36553 27568 36740
rect 27526 36544 27582 36553
rect 27526 36479 27582 36488
rect 27250 36408 27306 36417
rect 27250 36343 27306 36352
rect 27618 36272 27674 36281
rect 25872 36236 25924 36242
rect 27618 36207 27674 36216
rect 25872 36178 25924 36184
rect 25884 35873 25912 36178
rect 27632 36174 27660 36207
rect 27620 36168 27672 36174
rect 27620 36110 27672 36116
rect 28552 36038 28580 37431
rect 28644 37233 28672 41704
rect 28724 41686 28776 41692
rect 28828 41614 28856 42230
rect 29104 42158 29132 43862
rect 30564 43852 30616 43858
rect 30564 43794 30616 43800
rect 29552 43784 29604 43790
rect 29552 43726 29604 43732
rect 29920 43784 29972 43790
rect 29920 43726 29972 43732
rect 29564 43450 29592 43726
rect 29552 43444 29604 43450
rect 29552 43386 29604 43392
rect 29932 43382 29960 43726
rect 29920 43376 29972 43382
rect 29920 43318 29972 43324
rect 29932 43246 29960 43318
rect 29920 43240 29972 43246
rect 29920 43182 29972 43188
rect 30288 43240 30340 43246
rect 30288 43182 30340 43188
rect 30012 43104 30064 43110
rect 30012 43046 30064 43052
rect 30024 42906 30052 43046
rect 30012 42900 30064 42906
rect 30012 42842 30064 42848
rect 29460 42696 29512 42702
rect 29460 42638 29512 42644
rect 29092 42152 29144 42158
rect 29092 42094 29144 42100
rect 28724 41608 28776 41614
rect 28724 41550 28776 41556
rect 28816 41608 28868 41614
rect 28816 41550 28868 41556
rect 28736 39642 28764 41550
rect 29104 41414 29132 42094
rect 29472 41818 29500 42638
rect 29642 41984 29698 41993
rect 29642 41919 29698 41928
rect 29460 41812 29512 41818
rect 29460 41754 29512 41760
rect 29182 41712 29238 41721
rect 29182 41647 29184 41656
rect 29236 41647 29238 41656
rect 29184 41618 29236 41624
rect 29012 41386 29132 41414
rect 28908 41132 28960 41138
rect 28908 41074 28960 41080
rect 28724 39636 28776 39642
rect 28724 39578 28776 39584
rect 28920 39522 28948 41074
rect 29012 40594 29040 41386
rect 29472 40934 29500 41754
rect 29656 41750 29684 41919
rect 29644 41744 29696 41750
rect 29644 41686 29696 41692
rect 29828 41608 29880 41614
rect 29828 41550 29880 41556
rect 29460 40928 29512 40934
rect 29460 40870 29512 40876
rect 29840 40594 29868 41550
rect 30012 41132 30064 41138
rect 30012 41074 30064 41080
rect 30024 40934 30052 41074
rect 29920 40928 29972 40934
rect 29920 40870 29972 40876
rect 30012 40928 30064 40934
rect 30012 40870 30064 40876
rect 29932 40730 29960 40870
rect 29920 40724 29972 40730
rect 29920 40666 29972 40672
rect 29000 40588 29052 40594
rect 29000 40530 29052 40536
rect 29828 40588 29880 40594
rect 29828 40530 29880 40536
rect 29368 40384 29420 40390
rect 29368 40326 29420 40332
rect 29380 39642 29408 40326
rect 29840 40186 29868 40530
rect 29828 40180 29880 40186
rect 29828 40122 29880 40128
rect 29552 39976 29604 39982
rect 29552 39918 29604 39924
rect 29368 39636 29420 39642
rect 29368 39578 29420 39584
rect 28736 39506 28948 39522
rect 28724 39500 28948 39506
rect 28776 39494 28948 39500
rect 28724 39442 28776 39448
rect 28736 37262 28764 39442
rect 28816 39432 28868 39438
rect 28920 39420 28948 39494
rect 29000 39432 29052 39438
rect 28920 39392 29000 39420
rect 28816 39374 28868 39380
rect 29000 39374 29052 39380
rect 28828 38214 28856 39374
rect 29000 39296 29052 39302
rect 29000 39238 29052 39244
rect 29092 39296 29144 39302
rect 29092 39238 29144 39244
rect 29012 38826 29040 39238
rect 28908 38820 28960 38826
rect 28908 38762 28960 38768
rect 29000 38820 29052 38826
rect 29000 38762 29052 38768
rect 28816 38208 28868 38214
rect 28816 38150 28868 38156
rect 28828 37482 28856 38150
rect 28920 37942 28948 38762
rect 29104 38758 29132 39238
rect 29092 38752 29144 38758
rect 29092 38694 29144 38700
rect 29184 38752 29236 38758
rect 29184 38694 29236 38700
rect 29196 38486 29224 38694
rect 29564 38554 29592 39918
rect 30104 39432 30156 39438
rect 30104 39374 30156 39380
rect 30116 38962 30144 39374
rect 30300 38962 30328 43182
rect 30576 43110 30604 43794
rect 31036 43654 31064 44270
rect 31300 44192 31352 44198
rect 31300 44134 31352 44140
rect 31024 43648 31076 43654
rect 31024 43590 31076 43596
rect 30564 43104 30616 43110
rect 30564 43046 30616 43052
rect 30576 42906 30604 43046
rect 30564 42900 30616 42906
rect 30564 42842 30616 42848
rect 30656 42832 30708 42838
rect 30656 42774 30708 42780
rect 30472 42696 30524 42702
rect 30472 42638 30524 42644
rect 30380 42016 30432 42022
rect 30380 41958 30432 41964
rect 30392 41721 30420 41958
rect 30378 41712 30434 41721
rect 30378 41647 30434 41656
rect 30378 41576 30434 41585
rect 30378 41511 30434 41520
rect 30392 41478 30420 41511
rect 30380 41472 30432 41478
rect 30380 41414 30432 41420
rect 30380 41268 30432 41274
rect 30380 41210 30432 41216
rect 30392 41177 30420 41210
rect 30378 41168 30434 41177
rect 30378 41103 30434 41112
rect 30484 40934 30512 42638
rect 30668 42129 30696 42774
rect 31036 42770 31064 43590
rect 31312 43194 31340 44134
rect 32968 43994 32996 44474
rect 33416 44328 33468 44334
rect 33416 44270 33468 44276
rect 34336 44328 34388 44334
rect 34336 44270 34388 44276
rect 33324 44260 33376 44266
rect 33324 44202 33376 44208
rect 33232 44192 33284 44198
rect 33232 44134 33284 44140
rect 32956 43988 33008 43994
rect 32956 43930 33008 43936
rect 32220 43920 32272 43926
rect 32220 43862 32272 43868
rect 31760 43648 31812 43654
rect 31760 43590 31812 43596
rect 31772 43314 31800 43590
rect 31760 43308 31812 43314
rect 31220 43178 31340 43194
rect 31208 43172 31340 43178
rect 31260 43166 31340 43172
rect 31588 43268 31760 43296
rect 31208 43114 31260 43120
rect 31024 42764 31076 42770
rect 31024 42706 31076 42712
rect 30654 42120 30710 42129
rect 30654 42055 30710 42064
rect 30654 41984 30710 41993
rect 30654 41919 30710 41928
rect 30668 41313 30696 41919
rect 30654 41304 30710 41313
rect 30654 41239 30710 41248
rect 30932 41132 30984 41138
rect 30932 41074 30984 41080
rect 30564 41064 30616 41070
rect 30564 41006 30616 41012
rect 30472 40928 30524 40934
rect 30472 40870 30524 40876
rect 30380 39568 30432 39574
rect 30380 39510 30432 39516
rect 30392 39137 30420 39510
rect 30378 39128 30434 39137
rect 30378 39063 30434 39072
rect 30484 38962 30512 40870
rect 30576 40390 30604 41006
rect 30840 40588 30892 40594
rect 30840 40530 30892 40536
rect 30564 40384 30616 40390
rect 30564 40326 30616 40332
rect 30656 40384 30708 40390
rect 30656 40326 30708 40332
rect 30104 38956 30156 38962
rect 30104 38898 30156 38904
rect 30288 38956 30340 38962
rect 30288 38898 30340 38904
rect 30472 38956 30524 38962
rect 30472 38898 30524 38904
rect 29920 38752 29972 38758
rect 29920 38694 29972 38700
rect 29932 38554 29960 38694
rect 29552 38548 29604 38554
rect 29552 38490 29604 38496
rect 29920 38548 29972 38554
rect 29920 38490 29972 38496
rect 29184 38480 29236 38486
rect 29184 38422 29236 38428
rect 28908 37936 28960 37942
rect 28908 37878 28960 37884
rect 30196 37732 30248 37738
rect 30196 37674 30248 37680
rect 28906 37496 28962 37505
rect 28828 37454 28906 37482
rect 30208 37466 30236 37674
rect 28906 37431 28908 37440
rect 28960 37431 28962 37440
rect 30196 37460 30248 37466
rect 28908 37402 28960 37408
rect 30196 37402 30248 37408
rect 28998 37360 29054 37369
rect 28998 37295 29054 37304
rect 28724 37256 28776 37262
rect 28630 37224 28686 37233
rect 28724 37198 28776 37204
rect 28630 37159 28686 37168
rect 29012 36922 29040 37295
rect 30300 37194 30328 38898
rect 30576 38808 30604 40326
rect 30668 40186 30696 40326
rect 30656 40180 30708 40186
rect 30656 40122 30708 40128
rect 30852 39438 30880 40530
rect 30840 39432 30892 39438
rect 30840 39374 30892 39380
rect 30656 38820 30708 38826
rect 30576 38780 30656 38808
rect 30656 38762 30708 38768
rect 30288 37188 30340 37194
rect 30288 37130 30340 37136
rect 29000 36916 29052 36922
rect 29000 36858 29052 36864
rect 29000 36440 29052 36446
rect 29000 36382 29052 36388
rect 28540 36032 28592 36038
rect 28540 35974 28592 35980
rect 23572 35838 23624 35844
rect 25502 35864 25558 35873
rect 23202 35799 23258 35808
rect 23020 35760 23072 35766
rect 20074 35728 20130 35737
rect 20074 35663 20130 35672
rect 21178 35728 21234 35737
rect 21178 35663 21234 35672
rect 22006 35728 22062 35737
rect 22006 35663 22062 35672
rect 22190 35728 22246 35737
rect 22190 35663 22246 35672
rect 23018 35728 23020 35737
rect 23584 35737 23612 35838
rect 25502 35799 25558 35808
rect 25870 35864 25926 35873
rect 29012 35834 29040 36382
rect 30288 36372 30340 36378
rect 30288 36314 30340 36320
rect 29092 36032 29144 36038
rect 29092 35974 29144 35980
rect 25870 35799 25926 35808
rect 29000 35828 29052 35834
rect 29000 35770 29052 35776
rect 29104 35766 29132 35974
rect 30012 35896 30064 35902
rect 30300 35873 30328 36314
rect 30668 36009 30696 38762
rect 30838 38584 30894 38593
rect 30838 38519 30894 38528
rect 30748 38344 30800 38350
rect 30748 38286 30800 38292
rect 30760 37466 30788 38286
rect 30852 37913 30880 38519
rect 30838 37904 30894 37913
rect 30838 37839 30894 37848
rect 30748 37460 30800 37466
rect 30748 37402 30800 37408
rect 30840 37460 30892 37466
rect 30840 37402 30892 37408
rect 30852 37346 30880 37402
rect 30760 37330 30880 37346
rect 30748 37324 30880 37330
rect 30800 37318 30880 37324
rect 30748 37266 30800 37272
rect 30944 36009 30972 41074
rect 31024 40928 31076 40934
rect 31024 40870 31076 40876
rect 31036 40730 31064 40870
rect 31024 40724 31076 40730
rect 31024 40666 31076 40672
rect 31116 40520 31168 40526
rect 31116 40462 31168 40468
rect 31024 39840 31076 39846
rect 31024 39782 31076 39788
rect 30654 36000 30710 36009
rect 30654 35935 30710 35944
rect 30930 36000 30986 36009
rect 30930 35935 30986 35944
rect 30012 35838 30064 35844
rect 30286 35864 30342 35873
rect 29092 35760 29144 35766
rect 23072 35728 23074 35737
rect 23018 35663 23074 35672
rect 23570 35728 23626 35737
rect 30024 35737 30052 35838
rect 30286 35799 30342 35808
rect 31036 35737 31064 39782
rect 31128 39030 31156 40462
rect 31116 39024 31168 39030
rect 31116 38966 31168 38972
rect 31220 38486 31248 43114
rect 31300 43104 31352 43110
rect 31300 43046 31352 43052
rect 31312 42770 31340 43046
rect 31300 42764 31352 42770
rect 31300 42706 31352 42712
rect 31312 40526 31340 42706
rect 31484 41064 31536 41070
rect 31484 41006 31536 41012
rect 31392 40928 31444 40934
rect 31392 40870 31444 40876
rect 31300 40520 31352 40526
rect 31300 40462 31352 40468
rect 31298 40216 31354 40225
rect 31298 40151 31354 40160
rect 31208 38480 31260 38486
rect 31208 38422 31260 38428
rect 31208 37936 31260 37942
rect 31208 37878 31260 37884
rect 31220 37670 31248 37878
rect 31208 37664 31260 37670
rect 31208 37606 31260 37612
rect 31312 36922 31340 40151
rect 31404 39001 31432 40870
rect 31496 40186 31524 41006
rect 31484 40180 31536 40186
rect 31484 40122 31536 40128
rect 31496 39642 31524 40122
rect 31484 39636 31536 39642
rect 31484 39578 31536 39584
rect 31588 39506 31616 43268
rect 31760 43250 31812 43256
rect 32036 43172 32088 43178
rect 32036 43114 32088 43120
rect 31760 42900 31812 42906
rect 31760 42842 31812 42848
rect 31772 42158 31800 42842
rect 31852 42696 31904 42702
rect 31852 42638 31904 42644
rect 31760 42152 31812 42158
rect 31760 42094 31812 42100
rect 31772 41614 31800 42094
rect 31864 42022 31892 42638
rect 32048 42634 32076 43114
rect 32036 42628 32088 42634
rect 32036 42570 32088 42576
rect 32232 42226 32260 43862
rect 33244 43790 33272 44134
rect 33336 43926 33364 44202
rect 33428 43994 33456 44270
rect 33416 43988 33468 43994
rect 33416 43930 33468 43936
rect 33324 43920 33376 43926
rect 33324 43862 33376 43868
rect 33232 43784 33284 43790
rect 33232 43726 33284 43732
rect 34152 43784 34204 43790
rect 34152 43726 34204 43732
rect 34164 43450 34192 43726
rect 34152 43444 34204 43450
rect 34152 43386 34204 43392
rect 34242 43344 34298 43353
rect 33324 43308 33376 43314
rect 34242 43279 34298 43288
rect 33324 43250 33376 43256
rect 32496 43172 32548 43178
rect 32496 43114 32548 43120
rect 32508 42906 32536 43114
rect 32496 42900 32548 42906
rect 32496 42842 32548 42848
rect 32588 42900 32640 42906
rect 32588 42842 32640 42848
rect 33048 42900 33100 42906
rect 33048 42842 33100 42848
rect 32600 42786 32628 42842
rect 32312 42764 32364 42770
rect 32416 42758 32628 42786
rect 32416 42752 32444 42758
rect 32364 42724 32444 42752
rect 32312 42706 32364 42712
rect 33060 42362 33088 42842
rect 33232 42696 33284 42702
rect 33232 42638 33284 42644
rect 33244 42362 33272 42638
rect 33048 42356 33100 42362
rect 33048 42298 33100 42304
rect 33232 42356 33284 42362
rect 33232 42298 33284 42304
rect 32128 42220 32180 42226
rect 32128 42162 32180 42168
rect 32220 42220 32272 42226
rect 33232 42220 33284 42226
rect 32220 42162 32272 42168
rect 33060 42180 33232 42208
rect 32034 42120 32090 42129
rect 32034 42055 32090 42064
rect 31852 42016 31904 42022
rect 31852 41958 31904 41964
rect 32048 41750 32076 42055
rect 32036 41744 32088 41750
rect 32036 41686 32088 41692
rect 31760 41608 31812 41614
rect 31760 41550 31812 41556
rect 31668 40588 31720 40594
rect 31668 40530 31720 40536
rect 31760 40588 31812 40594
rect 31760 40530 31812 40536
rect 31576 39500 31628 39506
rect 31576 39442 31628 39448
rect 31680 39386 31708 40530
rect 31496 39358 31708 39386
rect 31390 38992 31446 39001
rect 31390 38927 31446 38936
rect 31392 38480 31444 38486
rect 31392 38422 31444 38428
rect 31404 37874 31432 38422
rect 31496 37913 31524 39358
rect 31574 39264 31630 39273
rect 31574 39199 31630 39208
rect 31482 37904 31538 37913
rect 31392 37868 31444 37874
rect 31482 37839 31538 37848
rect 31392 37810 31444 37816
rect 31496 37262 31524 37839
rect 31484 37256 31536 37262
rect 31484 37198 31536 37204
rect 31300 36916 31352 36922
rect 31300 36858 31352 36864
rect 31588 35766 31616 39199
rect 31668 38888 31720 38894
rect 31668 38830 31720 38836
rect 31680 37670 31708 38830
rect 31772 37874 31800 40530
rect 31852 40044 31904 40050
rect 31852 39986 31904 39992
rect 31864 39953 31892 39986
rect 31850 39944 31906 39953
rect 31850 39879 31906 39888
rect 31944 38820 31996 38826
rect 31944 38762 31996 38768
rect 31956 38729 31984 38762
rect 32140 38729 32168 42162
rect 32232 41750 32260 42162
rect 32864 42084 32916 42090
rect 32864 42026 32916 42032
rect 32220 41744 32272 41750
rect 32220 41686 32272 41692
rect 32232 40730 32260 41686
rect 32876 41682 32904 42026
rect 32864 41676 32916 41682
rect 32864 41618 32916 41624
rect 32956 41676 33008 41682
rect 32956 41618 33008 41624
rect 32588 41608 32640 41614
rect 32588 41550 32640 41556
rect 32680 41608 32732 41614
rect 32680 41550 32732 41556
rect 32220 40724 32272 40730
rect 32220 40666 32272 40672
rect 32600 40050 32628 41550
rect 32588 40044 32640 40050
rect 32588 39986 32640 39992
rect 32600 39914 32628 39986
rect 32588 39908 32640 39914
rect 32588 39850 32640 39856
rect 32220 39432 32272 39438
rect 32220 39374 32272 39380
rect 32588 39432 32640 39438
rect 32692 39420 32720 41550
rect 32968 41274 32996 41618
rect 33060 41614 33088 42180
rect 33232 42162 33284 42168
rect 33232 42016 33284 42022
rect 33232 41958 33284 41964
rect 33244 41818 33272 41958
rect 33140 41812 33192 41818
rect 33140 41754 33192 41760
rect 33232 41812 33284 41818
rect 33232 41754 33284 41760
rect 33152 41614 33180 41754
rect 33048 41608 33100 41614
rect 33048 41550 33100 41556
rect 33140 41608 33192 41614
rect 33140 41550 33192 41556
rect 32956 41268 33008 41274
rect 32956 41210 33008 41216
rect 32772 40996 32824 41002
rect 32772 40938 32824 40944
rect 32784 40730 32812 40938
rect 32968 40934 32996 41210
rect 33336 41177 33364 43250
rect 33508 42764 33560 42770
rect 33508 42706 33560 42712
rect 34060 42764 34112 42770
rect 34060 42706 34112 42712
rect 33416 42628 33468 42634
rect 33416 42570 33468 42576
rect 33322 41168 33378 41177
rect 33232 41132 33284 41138
rect 33428 41138 33456 42570
rect 33520 42362 33548 42706
rect 33600 42696 33652 42702
rect 33600 42638 33652 42644
rect 33508 42356 33560 42362
rect 33508 42298 33560 42304
rect 33612 41818 33640 42638
rect 33784 42016 33836 42022
rect 33784 41958 33836 41964
rect 33600 41812 33652 41818
rect 33600 41754 33652 41760
rect 33322 41103 33378 41112
rect 33416 41132 33468 41138
rect 33232 41074 33284 41080
rect 33416 41074 33468 41080
rect 32956 40928 33008 40934
rect 32956 40870 33008 40876
rect 33048 40928 33100 40934
rect 33048 40870 33100 40876
rect 32772 40724 32824 40730
rect 32772 40666 32824 40672
rect 33060 40186 33088 40870
rect 33140 40588 33192 40594
rect 33140 40530 33192 40536
rect 33048 40180 33100 40186
rect 33048 40122 33100 40128
rect 33152 40066 33180 40530
rect 33244 40390 33272 41074
rect 33692 41064 33744 41070
rect 33692 41006 33744 41012
rect 33600 40928 33652 40934
rect 33600 40870 33652 40876
rect 33508 40452 33560 40458
rect 33508 40394 33560 40400
rect 33232 40384 33284 40390
rect 33232 40326 33284 40332
rect 33520 40118 33548 40394
rect 32968 40038 33180 40066
rect 33508 40112 33560 40118
rect 33508 40054 33560 40060
rect 32968 39914 32996 40038
rect 32956 39908 33008 39914
rect 32956 39850 33008 39856
rect 32968 39506 32996 39850
rect 33612 39642 33640 40870
rect 33704 40730 33732 41006
rect 33796 41002 33824 41958
rect 34072 41614 34100 42706
rect 34256 41818 34284 43279
rect 34348 42906 34376 44270
rect 34428 44192 34480 44198
rect 34428 44134 34480 44140
rect 34520 44192 34572 44198
rect 34520 44134 34572 44140
rect 34440 43450 34468 44134
rect 34428 43444 34480 43450
rect 34428 43386 34480 43392
rect 34532 43246 34560 44134
rect 34520 43240 34572 43246
rect 34520 43182 34572 43188
rect 34428 43172 34480 43178
rect 34428 43114 34480 43120
rect 34336 42900 34388 42906
rect 34336 42842 34388 42848
rect 34440 42226 34468 43114
rect 34428 42220 34480 42226
rect 34428 42162 34480 42168
rect 34244 41812 34296 41818
rect 34244 41754 34296 41760
rect 34152 41676 34204 41682
rect 34152 41618 34204 41624
rect 34060 41608 34112 41614
rect 34060 41550 34112 41556
rect 34164 41138 34192 41618
rect 34152 41132 34204 41138
rect 34152 41074 34204 41080
rect 33784 40996 33836 41002
rect 33784 40938 33836 40944
rect 33692 40724 33744 40730
rect 33692 40666 33744 40672
rect 33704 39642 33732 40666
rect 33796 39914 33824 40938
rect 33968 40928 34020 40934
rect 33968 40870 34020 40876
rect 33980 40730 34008 40870
rect 33968 40724 34020 40730
rect 33968 40666 34020 40672
rect 34164 40526 34192 41074
rect 34426 40624 34482 40633
rect 34426 40559 34482 40568
rect 34060 40520 34112 40526
rect 34060 40462 34112 40468
rect 34152 40520 34204 40526
rect 34152 40462 34204 40468
rect 34072 40186 34100 40462
rect 34152 40384 34204 40390
rect 34152 40326 34204 40332
rect 34060 40180 34112 40186
rect 34060 40122 34112 40128
rect 33784 39908 33836 39914
rect 33784 39850 33836 39856
rect 33232 39636 33284 39642
rect 33232 39578 33284 39584
rect 33600 39636 33652 39642
rect 33600 39578 33652 39584
rect 33692 39636 33744 39642
rect 33692 39578 33744 39584
rect 32956 39500 33008 39506
rect 32956 39442 33008 39448
rect 32640 39392 32720 39420
rect 32588 39374 32640 39380
rect 32232 38962 32260 39374
rect 33244 39370 33272 39578
rect 33416 39500 33468 39506
rect 33416 39442 33468 39448
rect 33232 39364 33284 39370
rect 33232 39306 33284 39312
rect 32404 39296 32456 39302
rect 32404 39238 32456 39244
rect 32220 38956 32272 38962
rect 32220 38898 32272 38904
rect 32416 38894 32444 39238
rect 33046 38992 33102 39001
rect 33046 38927 33102 38936
rect 32404 38888 32456 38894
rect 32404 38830 32456 38836
rect 31942 38720 31998 38729
rect 31942 38655 31998 38664
rect 32126 38720 32182 38729
rect 32126 38655 32182 38664
rect 32956 38412 33008 38418
rect 32956 38354 33008 38360
rect 32968 38214 32996 38354
rect 32956 38208 33008 38214
rect 32956 38150 33008 38156
rect 32036 38004 32088 38010
rect 32036 37946 32088 37952
rect 31760 37868 31812 37874
rect 31760 37810 31812 37816
rect 32048 37670 32076 37946
rect 32312 37868 32364 37874
rect 32312 37810 32364 37816
rect 32220 37732 32272 37738
rect 32324 37720 32352 37810
rect 32272 37692 32352 37720
rect 32404 37732 32456 37738
rect 32220 37674 32272 37680
rect 32404 37674 32456 37680
rect 31668 37664 31720 37670
rect 31668 37606 31720 37612
rect 32036 37664 32088 37670
rect 32036 37606 32088 37612
rect 31680 37330 31708 37606
rect 32310 37496 32366 37505
rect 32416 37466 32444 37674
rect 32310 37431 32312 37440
rect 32364 37431 32366 37440
rect 32404 37460 32456 37466
rect 32312 37402 32364 37408
rect 32404 37402 32456 37408
rect 31668 37324 31720 37330
rect 31668 37266 31720 37272
rect 31680 35873 31708 37266
rect 33060 36378 33088 38927
rect 33232 38820 33284 38826
rect 33232 38762 33284 38768
rect 33244 38654 33272 38762
rect 33244 38626 33364 38654
rect 33140 38548 33192 38554
rect 33140 38490 33192 38496
rect 33152 38185 33180 38490
rect 33230 38448 33286 38457
rect 33230 38383 33232 38392
rect 33284 38383 33286 38392
rect 33232 38354 33284 38360
rect 33232 38208 33284 38214
rect 33138 38176 33194 38185
rect 33232 38150 33284 38156
rect 33138 38111 33194 38120
rect 33244 37777 33272 38150
rect 33230 37768 33286 37777
rect 33230 37703 33286 37712
rect 33138 37496 33194 37505
rect 33138 37431 33194 37440
rect 33152 37262 33180 37431
rect 33336 37398 33364 38626
rect 33324 37392 33376 37398
rect 33324 37334 33376 37340
rect 33140 37256 33192 37262
rect 33140 37198 33192 37204
rect 33048 36372 33100 36378
rect 33048 36314 33100 36320
rect 33428 36145 33456 39442
rect 33508 39296 33560 39302
rect 33508 39238 33560 39244
rect 33520 38826 33548 39238
rect 33600 39024 33652 39030
rect 33600 38966 33652 38972
rect 33508 38820 33560 38826
rect 33508 38762 33560 38768
rect 33520 37398 33548 38762
rect 33612 38729 33640 38966
rect 33968 38888 34020 38894
rect 33968 38830 34020 38836
rect 33784 38820 33836 38826
rect 33784 38762 33836 38768
rect 33598 38720 33654 38729
rect 33598 38655 33654 38664
rect 33690 38176 33746 38185
rect 33690 38111 33746 38120
rect 33704 38010 33732 38111
rect 33692 38004 33744 38010
rect 33692 37946 33744 37952
rect 33796 37874 33824 38762
rect 33876 38480 33928 38486
rect 33876 38422 33928 38428
rect 33784 37868 33836 37874
rect 33784 37810 33836 37816
rect 33690 37768 33746 37777
rect 33796 37754 33824 37810
rect 33746 37726 33824 37754
rect 33888 37738 33916 38422
rect 33980 38010 34008 38830
rect 33968 38004 34020 38010
rect 33968 37946 34020 37952
rect 33980 37806 34008 37946
rect 33968 37800 34020 37806
rect 33968 37742 34020 37748
rect 33876 37732 33928 37738
rect 33690 37703 33746 37712
rect 33508 37392 33560 37398
rect 33508 37334 33560 37340
rect 33600 37324 33652 37330
rect 33704 37312 33732 37703
rect 33876 37674 33928 37680
rect 33652 37284 33732 37312
rect 33600 37266 33652 37272
rect 33414 36136 33470 36145
rect 33414 36071 33470 36080
rect 34164 35873 34192 40326
rect 34440 39817 34468 40559
rect 34520 40112 34572 40118
rect 34520 40054 34572 40060
rect 34426 39808 34482 39817
rect 34426 39743 34482 39752
rect 34532 39574 34560 40054
rect 34624 39642 34652 45047
rect 39396 45008 39448 45014
rect 39396 44950 39448 44956
rect 35164 44396 35216 44402
rect 35164 44338 35216 44344
rect 38292 44396 38344 44402
rect 38292 44338 38344 44344
rect 35072 43648 35124 43654
rect 35072 43590 35124 43596
rect 34796 43104 34848 43110
rect 34796 43046 34848 43052
rect 34808 42906 34836 43046
rect 34796 42900 34848 42906
rect 34796 42842 34848 42848
rect 34980 42696 35032 42702
rect 34980 42638 35032 42644
rect 34888 41744 34940 41750
rect 34888 41686 34940 41692
rect 34794 41440 34850 41449
rect 34794 41375 34850 41384
rect 34808 41274 34836 41375
rect 34796 41268 34848 41274
rect 34796 41210 34848 41216
rect 34704 41200 34756 41206
rect 34704 41142 34756 41148
rect 34716 40089 34744 41142
rect 34808 40662 34836 41210
rect 34796 40656 34848 40662
rect 34796 40598 34848 40604
rect 34900 40458 34928 41686
rect 34888 40452 34940 40458
rect 34888 40394 34940 40400
rect 34702 40080 34758 40089
rect 34702 40015 34758 40024
rect 34900 39982 34928 40394
rect 34992 40118 35020 42638
rect 35084 42158 35112 43590
rect 35176 43314 35204 44338
rect 35256 44328 35308 44334
rect 35256 44270 35308 44276
rect 36728 44328 36780 44334
rect 36728 44270 36780 44276
rect 35268 43926 35296 44270
rect 35532 44192 35584 44198
rect 35532 44134 35584 44140
rect 35808 44192 35860 44198
rect 35808 44134 35860 44140
rect 36544 44192 36596 44198
rect 36544 44134 36596 44140
rect 35256 43920 35308 43926
rect 35256 43862 35308 43868
rect 35268 43654 35296 43862
rect 35440 43852 35492 43858
rect 35440 43794 35492 43800
rect 35348 43784 35400 43790
rect 35348 43726 35400 43732
rect 35256 43648 35308 43654
rect 35256 43590 35308 43596
rect 35164 43308 35216 43314
rect 35164 43250 35216 43256
rect 35072 42152 35124 42158
rect 35072 42094 35124 42100
rect 35176 41414 35204 43250
rect 35268 43246 35296 43590
rect 35256 43240 35308 43246
rect 35256 43182 35308 43188
rect 35360 43110 35388 43726
rect 35452 43382 35480 43794
rect 35544 43654 35572 44134
rect 35820 43790 35848 44134
rect 36556 43994 36584 44134
rect 36740 43994 36768 44270
rect 37740 44260 37792 44266
rect 37740 44202 37792 44208
rect 36544 43988 36596 43994
rect 36544 43930 36596 43936
rect 36728 43988 36780 43994
rect 36728 43930 36780 43936
rect 36360 43920 36412 43926
rect 36360 43862 36412 43868
rect 35808 43784 35860 43790
rect 35808 43726 35860 43732
rect 35532 43648 35584 43654
rect 35532 43590 35584 43596
rect 35440 43376 35492 43382
rect 35440 43318 35492 43324
rect 35348 43104 35400 43110
rect 35348 43046 35400 43052
rect 35360 42634 35388 43046
rect 35544 42702 35572 43590
rect 36372 43450 36400 43862
rect 36360 43444 36412 43450
rect 36360 43386 36412 43392
rect 36174 43072 36230 43081
rect 36174 43007 36230 43016
rect 36188 42838 36216 43007
rect 36372 42838 36400 43386
rect 36740 42906 36768 43930
rect 37752 43926 37780 44202
rect 38200 44192 38252 44198
rect 38200 44134 38252 44140
rect 38212 43926 38240 44134
rect 37740 43920 37792 43926
rect 37740 43862 37792 43868
rect 38200 43920 38252 43926
rect 38200 43862 38252 43868
rect 37752 43178 37780 43862
rect 38304 43314 38332 44338
rect 38844 44328 38896 44334
rect 38844 44270 38896 44276
rect 38476 43784 38528 43790
rect 38476 43726 38528 43732
rect 38292 43308 38344 43314
rect 38292 43250 38344 43256
rect 37740 43172 37792 43178
rect 37740 43114 37792 43120
rect 37924 43172 37976 43178
rect 37924 43114 37976 43120
rect 36728 42900 36780 42906
rect 36728 42842 36780 42848
rect 36176 42832 36228 42838
rect 36176 42774 36228 42780
rect 36360 42832 36412 42838
rect 36360 42774 36412 42780
rect 35532 42696 35584 42702
rect 35532 42638 35584 42644
rect 35348 42628 35400 42634
rect 35348 42570 35400 42576
rect 35360 42294 35388 42570
rect 36188 42362 36216 42774
rect 36636 42764 36688 42770
rect 36636 42706 36688 42712
rect 36452 42560 36504 42566
rect 36452 42502 36504 42508
rect 36464 42362 36492 42502
rect 36176 42356 36228 42362
rect 36176 42298 36228 42304
rect 36452 42356 36504 42362
rect 36452 42298 36504 42304
rect 35348 42288 35400 42294
rect 35348 42230 35400 42236
rect 35898 42256 35954 42265
rect 35898 42191 35954 42200
rect 35624 42152 35676 42158
rect 35624 42094 35676 42100
rect 35176 41386 35480 41414
rect 34980 40112 35032 40118
rect 34980 40054 35032 40060
rect 34888 39976 34940 39982
rect 34808 39936 34888 39964
rect 34612 39636 34664 39642
rect 34612 39578 34664 39584
rect 34520 39568 34572 39574
rect 34520 39510 34572 39516
rect 34704 38752 34756 38758
rect 34704 38694 34756 38700
rect 34242 37904 34298 37913
rect 34716 37874 34744 38694
rect 34242 37839 34244 37848
rect 34296 37839 34298 37848
rect 34704 37868 34756 37874
rect 34244 37810 34296 37816
rect 34704 37810 34756 37816
rect 34702 37768 34758 37777
rect 34702 37703 34758 37712
rect 34716 37670 34744 37703
rect 34704 37664 34756 37670
rect 34704 37606 34756 37612
rect 34808 37330 34836 39936
rect 34888 39918 34940 39924
rect 34992 39930 35020 40054
rect 34992 39902 35112 39930
rect 34888 38752 34940 38758
rect 34888 38694 34940 38700
rect 34900 38554 34928 38694
rect 34978 38584 35034 38593
rect 34888 38548 34940 38554
rect 34978 38519 35034 38528
rect 34888 38490 34940 38496
rect 34888 38412 34940 38418
rect 34992 38400 35020 38519
rect 34940 38372 35020 38400
rect 34888 38354 34940 38360
rect 34888 38276 34940 38282
rect 34888 38218 34940 38224
rect 34900 37670 34928 38218
rect 34980 37868 35032 37874
rect 34980 37810 35032 37816
rect 34888 37664 34940 37670
rect 34888 37606 34940 37612
rect 34992 37398 35020 37810
rect 34980 37392 35032 37398
rect 34980 37334 35032 37340
rect 34796 37324 34848 37330
rect 34796 37266 34848 37272
rect 35084 37262 35112 39902
rect 35256 39636 35308 39642
rect 35256 39578 35308 39584
rect 35164 38344 35216 38350
rect 35164 38286 35216 38292
rect 35176 37874 35204 38286
rect 35164 37868 35216 37874
rect 35164 37810 35216 37816
rect 35268 37806 35296 39578
rect 35452 38350 35480 41386
rect 35636 41138 35664 42094
rect 35912 42090 35940 42191
rect 35900 42084 35952 42090
rect 35900 42026 35952 42032
rect 36084 42084 36136 42090
rect 36084 42026 36136 42032
rect 35992 41608 36044 41614
rect 35992 41550 36044 41556
rect 36004 41478 36032 41550
rect 35808 41472 35860 41478
rect 35808 41414 35860 41420
rect 35992 41472 36044 41478
rect 35992 41414 36044 41420
rect 35624 41132 35676 41138
rect 35624 41074 35676 41080
rect 35636 39914 35664 41074
rect 35820 40934 35848 41414
rect 35808 40928 35860 40934
rect 35808 40870 35860 40876
rect 35806 39944 35862 39953
rect 35624 39908 35676 39914
rect 35806 39879 35862 39888
rect 35624 39850 35676 39856
rect 35636 39370 35664 39850
rect 35624 39364 35676 39370
rect 35624 39306 35676 39312
rect 35636 38962 35664 39306
rect 35624 38956 35676 38962
rect 35624 38898 35676 38904
rect 35636 38593 35664 38898
rect 35622 38584 35678 38593
rect 35622 38519 35678 38528
rect 35440 38344 35492 38350
rect 35440 38286 35492 38292
rect 35716 38344 35768 38350
rect 35716 38286 35768 38292
rect 35256 37800 35308 37806
rect 35256 37742 35308 37748
rect 35164 37732 35216 37738
rect 35164 37674 35216 37680
rect 35348 37732 35400 37738
rect 35348 37674 35400 37680
rect 35176 37398 35204 37674
rect 35360 37641 35388 37674
rect 35346 37632 35402 37641
rect 35346 37567 35402 37576
rect 35452 37505 35480 38286
rect 35532 37868 35584 37874
rect 35532 37810 35584 37816
rect 35438 37496 35494 37505
rect 35438 37431 35494 37440
rect 35164 37392 35216 37398
rect 35164 37334 35216 37340
rect 35072 37256 35124 37262
rect 35072 37198 35124 37204
rect 34428 36644 34480 36650
rect 34428 36586 34480 36592
rect 34440 35873 34468 36586
rect 35544 36281 35572 37810
rect 35728 37262 35756 38286
rect 35820 37890 35848 39879
rect 36004 39642 36032 41414
rect 36096 41052 36124 42026
rect 36176 41812 36228 41818
rect 36176 41754 36228 41760
rect 36188 41698 36216 41754
rect 36188 41670 36492 41698
rect 36464 41614 36492 41670
rect 36452 41608 36504 41614
rect 36452 41550 36504 41556
rect 36544 41540 36596 41546
rect 36544 41482 36596 41488
rect 36176 41064 36228 41070
rect 36096 41024 36176 41052
rect 36096 40594 36124 41024
rect 36176 41006 36228 41012
rect 36176 40724 36228 40730
rect 36176 40666 36228 40672
rect 36084 40588 36136 40594
rect 36084 40530 36136 40536
rect 36096 39914 36124 40530
rect 36084 39908 36136 39914
rect 36084 39850 36136 39856
rect 35992 39636 36044 39642
rect 35992 39578 36044 39584
rect 35900 38820 35952 38826
rect 35900 38762 35952 38768
rect 35912 38554 35940 38762
rect 35900 38548 35952 38554
rect 35900 38490 35952 38496
rect 35820 37862 35940 37890
rect 35912 37806 35940 37862
rect 35900 37800 35952 37806
rect 35900 37742 35952 37748
rect 36188 37670 36216 40666
rect 36556 40662 36584 41482
rect 36648 41478 36676 42706
rect 36820 42696 36872 42702
rect 36820 42638 36872 42644
rect 37188 42696 37240 42702
rect 37188 42638 37240 42644
rect 36728 41676 36780 41682
rect 36728 41618 36780 41624
rect 36636 41472 36688 41478
rect 36636 41414 36688 41420
rect 36648 41206 36676 41414
rect 36636 41200 36688 41206
rect 36636 41142 36688 41148
rect 36740 41138 36768 41618
rect 36832 41614 36860 42638
rect 37094 42392 37150 42401
rect 37094 42327 37150 42336
rect 36820 41608 36872 41614
rect 36820 41550 36872 41556
rect 36912 41268 36964 41274
rect 36912 41210 36964 41216
rect 36728 41132 36780 41138
rect 36728 41074 36780 41080
rect 36740 41041 36768 41074
rect 36726 41032 36782 41041
rect 36726 40967 36782 40976
rect 36728 40724 36780 40730
rect 36728 40666 36780 40672
rect 36544 40656 36596 40662
rect 36544 40598 36596 40604
rect 36634 39672 36690 39681
rect 36634 39607 36690 39616
rect 36648 39574 36676 39607
rect 36636 39568 36688 39574
rect 36636 39510 36688 39516
rect 36740 39506 36768 40666
rect 36544 39500 36596 39506
rect 36544 39442 36596 39448
rect 36728 39500 36780 39506
rect 36728 39442 36780 39448
rect 36268 38480 36320 38486
rect 36268 38422 36320 38428
rect 36280 38010 36308 38422
rect 36268 38004 36320 38010
rect 36268 37946 36320 37952
rect 36452 37936 36504 37942
rect 36452 37878 36504 37884
rect 36176 37664 36228 37670
rect 36176 37606 36228 37612
rect 36464 37466 36492 37878
rect 36452 37460 36504 37466
rect 36452 37402 36504 37408
rect 35716 37256 35768 37262
rect 35716 37198 35768 37204
rect 35716 36916 35768 36922
rect 35716 36858 35768 36864
rect 35530 36272 35586 36281
rect 35530 36207 35586 36216
rect 31666 35864 31722 35873
rect 34150 35864 34206 35873
rect 31666 35799 31722 35808
rect 33140 35828 33192 35834
rect 34150 35799 34206 35808
rect 34426 35864 34482 35873
rect 35728 35834 35756 36858
rect 36556 36553 36584 39442
rect 36740 39370 36768 39442
rect 36728 39364 36780 39370
rect 36728 39306 36780 39312
rect 36726 39264 36782 39273
rect 36726 39199 36782 39208
rect 36740 37398 36768 39199
rect 36820 38752 36872 38758
rect 36820 38694 36872 38700
rect 36832 38554 36860 38694
rect 36820 38548 36872 38554
rect 36820 38490 36872 38496
rect 36832 37466 36860 38490
rect 36924 38010 36952 41210
rect 37004 40928 37056 40934
rect 37004 40870 37056 40876
rect 37016 39574 37044 40870
rect 37108 40390 37136 42327
rect 37200 42022 37228 42638
rect 37832 42628 37884 42634
rect 37832 42570 37884 42576
rect 37464 42560 37516 42566
rect 37464 42502 37516 42508
rect 37476 42226 37504 42502
rect 37464 42220 37516 42226
rect 37464 42162 37516 42168
rect 37740 42152 37792 42158
rect 37740 42094 37792 42100
rect 37188 42016 37240 42022
rect 37188 41958 37240 41964
rect 37200 41818 37228 41958
rect 37188 41812 37240 41818
rect 37188 41754 37240 41760
rect 37372 41608 37424 41614
rect 37372 41550 37424 41556
rect 37384 41414 37412 41550
rect 37292 41386 37412 41414
rect 37096 40384 37148 40390
rect 37096 40326 37148 40332
rect 37292 40050 37320 41386
rect 37648 41064 37700 41070
rect 37648 41006 37700 41012
rect 37372 40452 37424 40458
rect 37372 40394 37424 40400
rect 37384 40050 37412 40394
rect 37464 40180 37516 40186
rect 37464 40122 37516 40128
rect 37280 40044 37332 40050
rect 37280 39986 37332 39992
rect 37372 40044 37424 40050
rect 37372 39986 37424 39992
rect 37004 39568 37056 39574
rect 37004 39510 37056 39516
rect 37292 38894 37320 39986
rect 37476 39438 37504 40122
rect 37372 39432 37424 39438
rect 37372 39374 37424 39380
rect 37464 39432 37516 39438
rect 37464 39374 37516 39380
rect 37384 38962 37412 39374
rect 37464 39296 37516 39302
rect 37464 39238 37516 39244
rect 37556 39296 37608 39302
rect 37556 39238 37608 39244
rect 37372 38956 37424 38962
rect 37372 38898 37424 38904
rect 37280 38888 37332 38894
rect 37280 38830 37332 38836
rect 37476 38826 37504 39238
rect 37568 39030 37596 39238
rect 37660 39030 37688 41006
rect 37752 40458 37780 42094
rect 37844 40934 37872 42570
rect 37832 40928 37884 40934
rect 37832 40870 37884 40876
rect 37936 40730 37964 43114
rect 38108 42764 38160 42770
rect 38108 42706 38160 42712
rect 38120 41138 38148 42706
rect 38200 42560 38252 42566
rect 38200 42502 38252 42508
rect 38304 42514 38332 43250
rect 38384 43104 38436 43110
rect 38384 43046 38436 43052
rect 38396 42702 38424 43046
rect 38384 42696 38436 42702
rect 38384 42638 38436 42644
rect 38488 42634 38516 43726
rect 38568 43648 38620 43654
rect 38568 43590 38620 43596
rect 38580 43246 38608 43590
rect 38568 43240 38620 43246
rect 38568 43182 38620 43188
rect 38856 43178 38884 44270
rect 39304 44260 39356 44266
rect 39304 44202 39356 44208
rect 38844 43172 38896 43178
rect 38844 43114 38896 43120
rect 39316 43110 39344 44202
rect 39408 43994 39436 44950
rect 49998 44636 50306 44645
rect 49998 44634 50004 44636
rect 50060 44634 50084 44636
rect 50140 44634 50164 44636
rect 50220 44634 50244 44636
rect 50300 44634 50306 44636
rect 50060 44582 50062 44634
rect 50242 44582 50244 44634
rect 49998 44580 50004 44582
rect 50060 44580 50084 44582
rect 50140 44580 50164 44582
rect 50220 44580 50244 44582
rect 50300 44580 50306 44582
rect 49998 44571 50306 44580
rect 43444 44464 43496 44470
rect 43444 44406 43496 44412
rect 47400 44464 47452 44470
rect 47400 44406 47452 44412
rect 41420 44396 41472 44402
rect 41420 44338 41472 44344
rect 39948 44328 40000 44334
rect 39948 44270 40000 44276
rect 40316 44328 40368 44334
rect 40316 44270 40368 44276
rect 41236 44328 41288 44334
rect 41236 44270 41288 44276
rect 39488 44192 39540 44198
rect 39488 44134 39540 44140
rect 39396 43988 39448 43994
rect 39396 43930 39448 43936
rect 39408 43382 39436 43930
rect 39396 43376 39448 43382
rect 39396 43318 39448 43324
rect 39396 43172 39448 43178
rect 39396 43114 39448 43120
rect 39304 43104 39356 43110
rect 39304 43046 39356 43052
rect 38752 42696 38804 42702
rect 38752 42638 38804 42644
rect 38476 42628 38528 42634
rect 38476 42570 38528 42576
rect 38212 42158 38240 42502
rect 38304 42486 38424 42514
rect 38396 42226 38424 42486
rect 38384 42220 38436 42226
rect 38384 42162 38436 42168
rect 38200 42152 38252 42158
rect 38200 42094 38252 42100
rect 38396 41750 38424 42162
rect 38384 41744 38436 41750
rect 38384 41686 38436 41692
rect 38488 41682 38516 42570
rect 38476 41676 38528 41682
rect 38476 41618 38528 41624
rect 38488 41414 38516 41618
rect 38488 41386 38700 41414
rect 38108 41132 38160 41138
rect 38108 41074 38160 41080
rect 38476 41064 38528 41070
rect 38476 41006 38528 41012
rect 38108 40928 38160 40934
rect 38108 40870 38160 40876
rect 37924 40724 37976 40730
rect 37924 40666 37976 40672
rect 37740 40452 37792 40458
rect 37740 40394 37792 40400
rect 38120 40186 38148 40870
rect 38488 40662 38516 41006
rect 38476 40656 38528 40662
rect 38476 40598 38528 40604
rect 38108 40180 38160 40186
rect 38108 40122 38160 40128
rect 38108 39908 38160 39914
rect 38108 39850 38160 39856
rect 38120 39506 38148 39850
rect 38108 39500 38160 39506
rect 38108 39442 38160 39448
rect 37556 39024 37608 39030
rect 37556 38966 37608 38972
rect 37648 39024 37700 39030
rect 37648 38966 37700 38972
rect 37740 39024 37792 39030
rect 37740 38966 37792 38972
rect 37188 38820 37240 38826
rect 37188 38762 37240 38768
rect 37464 38820 37516 38826
rect 37464 38762 37516 38768
rect 37200 38282 37228 38762
rect 37372 38752 37424 38758
rect 37372 38694 37424 38700
rect 37384 38418 37412 38694
rect 37372 38412 37424 38418
rect 37372 38354 37424 38360
rect 37188 38276 37240 38282
rect 37188 38218 37240 38224
rect 37752 38162 37780 38966
rect 38292 38888 38344 38894
rect 38292 38830 38344 38836
rect 38304 38554 38332 38830
rect 38292 38548 38344 38554
rect 38292 38490 38344 38496
rect 37200 38134 37780 38162
rect 36912 38004 36964 38010
rect 36912 37946 36964 37952
rect 37004 38004 37056 38010
rect 37004 37946 37056 37952
rect 37016 37738 37044 37946
rect 37004 37732 37056 37738
rect 37004 37674 37056 37680
rect 36820 37460 36872 37466
rect 36820 37402 36872 37408
rect 36728 37392 36780 37398
rect 36728 37334 36780 37340
rect 37200 37233 37228 38134
rect 38304 37806 38332 38490
rect 37740 37800 37792 37806
rect 37740 37742 37792 37748
rect 38292 37800 38344 37806
rect 38292 37742 38344 37748
rect 37280 37664 37332 37670
rect 37280 37606 37332 37612
rect 37186 37224 37242 37233
rect 37186 37159 37242 37168
rect 37292 36650 37320 37606
rect 37752 36825 37780 37742
rect 38488 37262 38516 40598
rect 38672 40050 38700 41386
rect 38660 40044 38712 40050
rect 38660 39986 38712 39992
rect 38764 39681 38792 42638
rect 38844 42560 38896 42566
rect 38844 42502 38896 42508
rect 38856 41750 38884 42502
rect 39120 41812 39172 41818
rect 39120 41754 39172 41760
rect 38844 41744 38896 41750
rect 38844 41686 38896 41692
rect 38936 41472 38988 41478
rect 38936 41414 38988 41420
rect 38842 40216 38898 40225
rect 38842 40151 38898 40160
rect 38750 39672 38806 39681
rect 38568 39636 38620 39642
rect 38750 39607 38806 39616
rect 38568 39578 38620 39584
rect 38580 39438 38608 39578
rect 38568 39432 38620 39438
rect 38568 39374 38620 39380
rect 38764 39302 38792 39607
rect 38752 39296 38804 39302
rect 38752 39238 38804 39244
rect 38476 37256 38528 37262
rect 38476 37198 38528 37204
rect 38660 37120 38712 37126
rect 38660 37062 38712 37068
rect 37738 36816 37794 36825
rect 37738 36751 37794 36760
rect 37280 36644 37332 36650
rect 37280 36586 37332 36592
rect 36542 36544 36598 36553
rect 36542 36479 36598 36488
rect 38672 36281 38700 37062
rect 38856 36718 38884 40151
rect 38948 39642 38976 41414
rect 38936 39636 38988 39642
rect 38936 39578 38988 39584
rect 39132 39438 39160 41754
rect 39212 40928 39264 40934
rect 39212 40870 39264 40876
rect 39120 39432 39172 39438
rect 39120 39374 39172 39380
rect 39224 39030 39252 40870
rect 39212 39024 39264 39030
rect 39212 38966 39264 38972
rect 39316 38842 39344 43046
rect 39408 40118 39436 43114
rect 39500 42906 39528 44134
rect 39580 43104 39632 43110
rect 39580 43046 39632 43052
rect 39488 42900 39540 42906
rect 39488 42842 39540 42848
rect 39592 42090 39620 43046
rect 39580 42084 39632 42090
rect 39580 42026 39632 42032
rect 39960 41682 39988 44270
rect 40132 43308 40184 43314
rect 40132 43250 40184 43256
rect 40040 42560 40092 42566
rect 40040 42502 40092 42508
rect 39948 41676 40000 41682
rect 39948 41618 40000 41624
rect 40052 41206 40080 42502
rect 40040 41200 40092 41206
rect 40040 41142 40092 41148
rect 39580 41132 39632 41138
rect 39580 41074 39632 41080
rect 39488 40928 39540 40934
rect 39488 40870 39540 40876
rect 39500 40662 39528 40870
rect 39488 40656 39540 40662
rect 39488 40598 39540 40604
rect 39396 40112 39448 40118
rect 39396 40054 39448 40060
rect 39396 39024 39448 39030
rect 39396 38966 39448 38972
rect 39224 38814 39344 38842
rect 39120 38752 39172 38758
rect 39120 38694 39172 38700
rect 39132 37806 39160 38694
rect 39224 38486 39252 38814
rect 39212 38480 39264 38486
rect 39212 38422 39264 38428
rect 39224 38350 39252 38422
rect 39212 38344 39264 38350
rect 39212 38286 39264 38292
rect 39304 38344 39356 38350
rect 39304 38286 39356 38292
rect 39120 37800 39172 37806
rect 39120 37742 39172 37748
rect 39316 37670 39344 38286
rect 39304 37664 39356 37670
rect 39304 37606 39356 37612
rect 39408 37097 39436 38966
rect 39488 38956 39540 38962
rect 39488 38898 39540 38904
rect 39500 37874 39528 38898
rect 39592 38894 39620 41074
rect 39672 40928 39724 40934
rect 39672 40870 39724 40876
rect 39684 40508 39712 40870
rect 39856 40520 39908 40526
rect 39684 40480 39856 40508
rect 39684 40186 39712 40480
rect 39856 40462 39908 40468
rect 40052 40390 40080 41142
rect 40144 41138 40172 43250
rect 40328 43246 40356 44270
rect 40868 44192 40920 44198
rect 40868 44134 40920 44140
rect 40316 43240 40368 43246
rect 40236 43200 40316 43228
rect 40236 41614 40264 43200
rect 40316 43182 40368 43188
rect 40408 43104 40460 43110
rect 40408 43046 40460 43052
rect 40420 42906 40448 43046
rect 40408 42900 40460 42906
rect 40408 42842 40460 42848
rect 40592 42696 40644 42702
rect 40592 42638 40644 42644
rect 40776 42696 40828 42702
rect 40776 42638 40828 42644
rect 40604 42566 40632 42638
rect 40592 42560 40644 42566
rect 40592 42502 40644 42508
rect 40788 42362 40816 42638
rect 40776 42356 40828 42362
rect 40776 42298 40828 42304
rect 40316 42220 40368 42226
rect 40316 42162 40368 42168
rect 40328 41750 40356 42162
rect 40316 41744 40368 41750
rect 40316 41686 40368 41692
rect 40500 41744 40552 41750
rect 40500 41686 40552 41692
rect 40224 41608 40276 41614
rect 40224 41550 40276 41556
rect 40512 41138 40540 41686
rect 40776 41540 40828 41546
rect 40880 41528 40908 44134
rect 41248 43994 41276 44270
rect 41432 44198 41460 44338
rect 43352 44328 43404 44334
rect 43352 44270 43404 44276
rect 41420 44192 41472 44198
rect 41420 44134 41472 44140
rect 42156 44192 42208 44198
rect 42156 44134 42208 44140
rect 42340 44192 42392 44198
rect 42340 44134 42392 44140
rect 42524 44192 42576 44198
rect 42524 44134 42576 44140
rect 41236 43988 41288 43994
rect 41236 43930 41288 43936
rect 40960 43784 41012 43790
rect 40960 43726 41012 43732
rect 41236 43784 41288 43790
rect 41236 43726 41288 43732
rect 40972 43450 41000 43726
rect 40960 43444 41012 43450
rect 40960 43386 41012 43392
rect 41248 43382 41276 43726
rect 41236 43376 41288 43382
rect 41236 43318 41288 43324
rect 41432 43314 41460 44134
rect 42168 43926 42196 44134
rect 42156 43920 42208 43926
rect 42156 43862 42208 43868
rect 41880 43784 41932 43790
rect 41880 43726 41932 43732
rect 41420 43308 41472 43314
rect 41420 43250 41472 43256
rect 41144 42900 41196 42906
rect 41144 42842 41196 42848
rect 40960 42084 41012 42090
rect 40960 42026 41012 42032
rect 40972 41682 41000 42026
rect 41156 42022 41184 42842
rect 41432 42770 41460 43250
rect 41788 43104 41840 43110
rect 41786 43072 41788 43081
rect 41840 43072 41842 43081
rect 41786 43007 41842 43016
rect 41420 42764 41472 42770
rect 41420 42706 41472 42712
rect 41788 42764 41840 42770
rect 41788 42706 41840 42712
rect 41420 42628 41472 42634
rect 41420 42570 41472 42576
rect 41432 42158 41460 42570
rect 41420 42152 41472 42158
rect 41420 42094 41472 42100
rect 41512 42084 41564 42090
rect 41512 42026 41564 42032
rect 41144 42016 41196 42022
rect 41144 41958 41196 41964
rect 40960 41676 41012 41682
rect 40960 41618 41012 41624
rect 40828 41500 40908 41528
rect 40776 41482 40828 41488
rect 40684 41472 40736 41478
rect 40684 41414 40736 41420
rect 40696 41313 40724 41414
rect 40682 41304 40738 41313
rect 40682 41239 40738 41248
rect 40132 41132 40184 41138
rect 40132 41074 40184 41080
rect 40500 41132 40552 41138
rect 40500 41074 40552 41080
rect 39948 40384 40000 40390
rect 39948 40326 40000 40332
rect 40040 40384 40092 40390
rect 40040 40326 40092 40332
rect 39672 40180 39724 40186
rect 39672 40122 39724 40128
rect 39764 39976 39816 39982
rect 39764 39918 39816 39924
rect 39776 38894 39804 39918
rect 39580 38888 39632 38894
rect 39580 38830 39632 38836
rect 39764 38888 39816 38894
rect 39764 38830 39816 38836
rect 39672 38480 39724 38486
rect 39672 38422 39724 38428
rect 39684 37913 39712 38422
rect 39776 38298 39804 38830
rect 39960 38434 39988 40326
rect 40144 40202 40172 41074
rect 40512 41002 40540 41074
rect 40500 40996 40552 41002
rect 40500 40938 40552 40944
rect 40512 40730 40540 40938
rect 40500 40724 40552 40730
rect 40500 40666 40552 40672
rect 40144 40174 40264 40202
rect 40040 39908 40092 39914
rect 40040 39850 40092 39856
rect 40052 38554 40080 39850
rect 40132 39296 40184 39302
rect 40132 39238 40184 39244
rect 40144 39030 40172 39238
rect 40132 39024 40184 39030
rect 40132 38966 40184 38972
rect 40132 38752 40184 38758
rect 40132 38694 40184 38700
rect 40040 38548 40092 38554
rect 40040 38490 40092 38496
rect 39960 38406 40080 38434
rect 39948 38344 40000 38350
rect 39776 38292 39948 38298
rect 39776 38286 40000 38292
rect 39776 38270 39988 38286
rect 39670 37904 39726 37913
rect 39488 37868 39540 37874
rect 39670 37839 39726 37848
rect 39488 37810 39540 37816
rect 40052 37244 40080 38406
rect 40144 37806 40172 38694
rect 40236 38486 40264 40174
rect 40408 39364 40460 39370
rect 40408 39306 40460 39312
rect 40420 39030 40448 39306
rect 40408 39024 40460 39030
rect 40408 38966 40460 38972
rect 40512 38962 40724 38978
rect 40500 38956 40736 38962
rect 40552 38950 40684 38956
rect 40500 38898 40552 38904
rect 40684 38898 40736 38904
rect 40500 38752 40552 38758
rect 40500 38694 40552 38700
rect 40224 38480 40276 38486
rect 40224 38422 40276 38428
rect 40512 37806 40540 38694
rect 40788 37874 40816 41482
rect 40972 40662 41000 41618
rect 41052 40928 41104 40934
rect 41052 40870 41104 40876
rect 41064 40730 41092 40870
rect 41052 40724 41104 40730
rect 41052 40666 41104 40672
rect 40960 40656 41012 40662
rect 40960 40598 41012 40604
rect 40972 39964 41000 40598
rect 41052 39976 41104 39982
rect 40972 39936 41052 39964
rect 40972 39574 41000 39936
rect 41052 39918 41104 39924
rect 41052 39840 41104 39846
rect 41050 39808 41052 39817
rect 41104 39808 41106 39817
rect 41050 39743 41106 39752
rect 40960 39568 41012 39574
rect 40960 39510 41012 39516
rect 40972 39114 41000 39510
rect 41156 39386 41184 41958
rect 41524 40730 41552 42026
rect 41800 41614 41828 42706
rect 41892 42702 41920 43726
rect 42352 43450 42380 44134
rect 42340 43444 42392 43450
rect 42340 43386 42392 43392
rect 41972 43172 42024 43178
rect 41972 43114 42024 43120
rect 41984 42906 42012 43114
rect 42536 42906 42564 44134
rect 43168 43784 43220 43790
rect 43168 43726 43220 43732
rect 43076 43240 43128 43246
rect 43180 43228 43208 43726
rect 43364 43382 43392 44270
rect 43456 43926 43484 44406
rect 44364 44396 44416 44402
rect 44364 44338 44416 44344
rect 46112 44396 46164 44402
rect 46112 44338 46164 44344
rect 44180 44328 44232 44334
rect 44180 44270 44232 44276
rect 43444 43920 43496 43926
rect 43444 43862 43496 43868
rect 43904 43852 43956 43858
rect 43904 43794 43956 43800
rect 43812 43648 43864 43654
rect 43812 43590 43864 43596
rect 43824 43450 43852 43590
rect 43812 43444 43864 43450
rect 43812 43386 43864 43392
rect 43352 43376 43404 43382
rect 43352 43318 43404 43324
rect 43128 43200 43208 43228
rect 43076 43182 43128 43188
rect 41972 42900 42024 42906
rect 41972 42842 42024 42848
rect 42524 42900 42576 42906
rect 42524 42842 42576 42848
rect 43180 42838 43208 43200
rect 43168 42832 43220 42838
rect 42812 42780 43168 42786
rect 42812 42774 43220 42780
rect 42812 42758 43208 42774
rect 41880 42696 41932 42702
rect 41880 42638 41932 42644
rect 42156 42696 42208 42702
rect 42156 42638 42208 42644
rect 42524 42696 42576 42702
rect 42524 42638 42576 42644
rect 41892 42090 41920 42638
rect 41880 42084 41932 42090
rect 41880 42026 41932 42032
rect 41788 41608 41840 41614
rect 41788 41550 41840 41556
rect 41696 41132 41748 41138
rect 41696 41074 41748 41080
rect 41512 40724 41564 40730
rect 41512 40666 41564 40672
rect 41708 40458 41736 41074
rect 41892 40526 41920 42026
rect 42168 41818 42196 42638
rect 42536 41818 42564 42638
rect 42156 41812 42208 41818
rect 42156 41754 42208 41760
rect 42524 41812 42576 41818
rect 42524 41754 42576 41760
rect 42524 41608 42576 41614
rect 42524 41550 42576 41556
rect 42248 41064 42300 41070
rect 42248 41006 42300 41012
rect 41970 40760 42026 40769
rect 42260 40730 42288 41006
rect 42536 40882 42564 41550
rect 42708 41472 42760 41478
rect 42708 41414 42760 41420
rect 42720 41256 42748 41414
rect 42628 41228 42748 41256
rect 42628 41002 42656 41228
rect 42812 41002 42840 42758
rect 43260 42560 43312 42566
rect 43260 42502 43312 42508
rect 43628 42560 43680 42566
rect 43628 42502 43680 42508
rect 43168 42084 43220 42090
rect 43168 42026 43220 42032
rect 43074 41848 43130 41857
rect 43074 41783 43130 41792
rect 42616 40996 42668 41002
rect 42616 40938 42668 40944
rect 42800 40996 42852 41002
rect 42800 40938 42852 40944
rect 42536 40854 42656 40882
rect 41970 40695 42026 40704
rect 42064 40724 42116 40730
rect 41984 40594 42012 40695
rect 42064 40666 42116 40672
rect 42248 40724 42300 40730
rect 42248 40666 42300 40672
rect 41972 40588 42024 40594
rect 41972 40530 42024 40536
rect 41880 40520 41932 40526
rect 41880 40462 41932 40468
rect 41696 40452 41748 40458
rect 41696 40394 41748 40400
rect 41420 40180 41472 40186
rect 41420 40122 41472 40128
rect 41432 40032 41460 40122
rect 41604 40112 41656 40118
rect 41604 40054 41656 40060
rect 41064 39358 41184 39386
rect 41340 40004 41460 40032
rect 41064 39302 41092 39358
rect 41052 39296 41104 39302
rect 41052 39238 41104 39244
rect 41234 39264 41290 39273
rect 41234 39199 41290 39208
rect 40972 39086 41092 39114
rect 40960 38956 41012 38962
rect 40960 38898 41012 38904
rect 40776 37868 40828 37874
rect 40776 37810 40828 37816
rect 40972 37806 41000 38898
rect 41064 38758 41092 39086
rect 41052 38752 41104 38758
rect 41052 38694 41104 38700
rect 41050 38584 41106 38593
rect 41248 38554 41276 39199
rect 41340 38962 41368 40004
rect 41616 39964 41644 40054
rect 41432 39936 41644 39964
rect 41432 39438 41460 39936
rect 41512 39840 41564 39846
rect 41512 39782 41564 39788
rect 41604 39840 41656 39846
rect 41604 39782 41656 39788
rect 41524 39574 41552 39782
rect 41512 39568 41564 39574
rect 41512 39510 41564 39516
rect 41420 39432 41472 39438
rect 41420 39374 41472 39380
rect 41328 38956 41380 38962
rect 41328 38898 41380 38904
rect 41050 38519 41106 38528
rect 41236 38548 41288 38554
rect 41064 38214 41092 38519
rect 41236 38490 41288 38496
rect 41144 38480 41196 38486
rect 41144 38422 41196 38428
rect 41052 38208 41104 38214
rect 41052 38150 41104 38156
rect 40132 37800 40184 37806
rect 40132 37742 40184 37748
rect 40500 37800 40552 37806
rect 40500 37742 40552 37748
rect 40960 37800 41012 37806
rect 40960 37742 41012 37748
rect 40132 37664 40184 37670
rect 40132 37606 40184 37612
rect 40144 37398 40172 37606
rect 40132 37392 40184 37398
rect 40132 37334 40184 37340
rect 41156 37312 41184 38422
rect 41236 38412 41288 38418
rect 41236 38354 41288 38360
rect 41328 38412 41380 38418
rect 41328 38354 41380 38360
rect 41248 38010 41276 38354
rect 41236 38004 41288 38010
rect 41236 37946 41288 37952
rect 41340 37913 41368 38354
rect 41326 37904 41382 37913
rect 41326 37839 41382 37848
rect 41340 37330 41368 37839
rect 41524 37806 41552 39510
rect 41616 39273 41644 39782
rect 41708 39386 41736 40394
rect 42076 40390 42104 40666
rect 42248 40588 42300 40594
rect 42248 40530 42300 40536
rect 42064 40384 42116 40390
rect 42064 40326 42116 40332
rect 42156 39976 42208 39982
rect 42156 39918 42208 39924
rect 41972 39840 42024 39846
rect 41972 39782 42024 39788
rect 41788 39432 41840 39438
rect 41708 39380 41788 39386
rect 41708 39374 41840 39380
rect 41880 39432 41932 39438
rect 41880 39374 41932 39380
rect 41708 39358 41828 39374
rect 41602 39264 41658 39273
rect 41602 39199 41658 39208
rect 41708 38282 41736 39358
rect 41788 39296 41840 39302
rect 41788 39238 41840 39244
rect 41800 38826 41828 39238
rect 41788 38820 41840 38826
rect 41788 38762 41840 38768
rect 41892 38350 41920 39374
rect 41984 39370 42012 39782
rect 42168 39370 42196 39918
rect 41972 39364 42024 39370
rect 41972 39306 42024 39312
rect 42156 39364 42208 39370
rect 42156 39306 42208 39312
rect 41880 38344 41932 38350
rect 41880 38286 41932 38292
rect 41970 38312 42026 38321
rect 41696 38276 41748 38282
rect 41970 38247 42026 38256
rect 41696 38218 41748 38224
rect 41512 37800 41564 37806
rect 41512 37742 41564 37748
rect 41604 37664 41656 37670
rect 41604 37606 41656 37612
rect 41616 37346 41644 37606
rect 41708 37466 41736 38218
rect 41984 38214 42012 38247
rect 41972 38208 42024 38214
rect 41972 38150 42024 38156
rect 41984 37806 42012 38150
rect 41972 37800 42024 37806
rect 41972 37742 42024 37748
rect 42168 37670 42196 39306
rect 42156 37664 42208 37670
rect 42156 37606 42208 37612
rect 41696 37460 41748 37466
rect 41696 37402 41748 37408
rect 41236 37324 41288 37330
rect 41156 37284 41236 37312
rect 41236 37266 41288 37272
rect 41328 37324 41380 37330
rect 41616 37318 41736 37346
rect 41328 37266 41380 37272
rect 40052 37216 40172 37244
rect 39394 37088 39450 37097
rect 39394 37023 39450 37032
rect 38844 36712 38896 36718
rect 38844 36654 38896 36660
rect 38658 36272 38714 36281
rect 38658 36207 38714 36216
rect 38658 36136 38714 36145
rect 38658 36071 38660 36080
rect 38712 36071 38714 36080
rect 38660 36042 38712 36048
rect 35806 36000 35862 36009
rect 35806 35935 35808 35944
rect 35860 35935 35862 35944
rect 35808 35906 35860 35912
rect 40144 35873 40172 37216
rect 41708 37126 41736 37318
rect 41696 37120 41748 37126
rect 41696 37062 41748 37068
rect 41708 36689 41736 37062
rect 42260 36922 42288 40530
rect 42432 39500 42484 39506
rect 42432 39442 42484 39448
rect 42340 39296 42392 39302
rect 42340 39238 42392 39244
rect 42352 39098 42380 39238
rect 42444 39098 42472 39442
rect 42628 39438 42656 40854
rect 42892 40656 42944 40662
rect 42892 40598 42944 40604
rect 42904 39658 42932 40598
rect 43088 40050 43116 41783
rect 43180 41614 43208 42026
rect 43168 41608 43220 41614
rect 43168 41550 43220 41556
rect 43272 41478 43300 42502
rect 43444 42084 43496 42090
rect 43444 42026 43496 42032
rect 43352 41812 43404 41818
rect 43352 41754 43404 41760
rect 43260 41472 43312 41478
rect 43260 41414 43312 41420
rect 43168 40996 43220 41002
rect 43168 40938 43220 40944
rect 43180 40662 43208 40938
rect 43168 40656 43220 40662
rect 43168 40598 43220 40604
rect 43364 40186 43392 41754
rect 43456 41274 43484 42026
rect 43536 41812 43588 41818
rect 43536 41754 43588 41760
rect 43548 41721 43576 41754
rect 43640 41750 43668 42502
rect 43916 42362 43944 43794
rect 44192 43722 44220 44270
rect 44180 43716 44232 43722
rect 44180 43658 44232 43664
rect 43996 43308 44048 43314
rect 43996 43250 44048 43256
rect 44088 43308 44140 43314
rect 44088 43250 44140 43256
rect 44008 42906 44036 43250
rect 43996 42900 44048 42906
rect 43996 42842 44048 42848
rect 44100 42770 44128 43250
rect 44270 43072 44326 43081
rect 44270 43007 44326 43016
rect 44088 42764 44140 42770
rect 44088 42706 44140 42712
rect 43904 42356 43956 42362
rect 43904 42298 43956 42304
rect 43916 41818 43944 42298
rect 44100 42226 44128 42706
rect 44180 42696 44232 42702
rect 44180 42638 44232 42644
rect 44088 42220 44140 42226
rect 44088 42162 44140 42168
rect 43812 41812 43864 41818
rect 43812 41754 43864 41760
rect 43904 41812 43956 41818
rect 43904 41754 43956 41760
rect 43628 41744 43680 41750
rect 43534 41712 43590 41721
rect 43628 41686 43680 41692
rect 43824 41682 43852 41754
rect 43534 41647 43590 41656
rect 43812 41676 43864 41682
rect 43812 41618 43864 41624
rect 43812 41472 43864 41478
rect 43812 41414 43864 41420
rect 43916 41414 43944 41754
rect 44100 41478 44128 42162
rect 44088 41472 44140 41478
rect 44088 41414 44140 41420
rect 44192 41414 44220 42638
rect 44284 42362 44312 43007
rect 44272 42356 44324 42362
rect 44272 42298 44324 42304
rect 44270 42120 44326 42129
rect 44270 42055 44272 42064
rect 44324 42055 44326 42064
rect 44272 42026 44324 42032
rect 43444 41268 43496 41274
rect 43444 41210 43496 41216
rect 43720 40384 43772 40390
rect 43720 40326 43772 40332
rect 43352 40180 43404 40186
rect 43352 40122 43404 40128
rect 43076 40044 43128 40050
rect 43076 39986 43128 39992
rect 43536 40044 43588 40050
rect 43536 39986 43588 39992
rect 43548 39846 43576 39986
rect 43732 39846 43760 40326
rect 43824 40118 43852 41414
rect 43916 41386 44036 41414
rect 44192 41386 44312 41414
rect 43902 41304 43958 41313
rect 43902 41239 43958 41248
rect 43812 40112 43864 40118
rect 43812 40054 43864 40060
rect 43536 39840 43588 39846
rect 43536 39782 43588 39788
rect 43720 39840 43772 39846
rect 43720 39782 43772 39788
rect 42904 39642 43024 39658
rect 42904 39636 43036 39642
rect 42904 39630 42984 39636
rect 42984 39578 43036 39584
rect 43444 39568 43496 39574
rect 43444 39510 43496 39516
rect 42708 39500 42760 39506
rect 42708 39442 42760 39448
rect 42616 39432 42668 39438
rect 42616 39374 42668 39380
rect 42340 39092 42392 39098
rect 42340 39034 42392 39040
rect 42432 39092 42484 39098
rect 42432 39034 42484 39040
rect 42524 38956 42576 38962
rect 42524 38898 42576 38904
rect 42536 38554 42564 38898
rect 42524 38548 42576 38554
rect 42524 38490 42576 38496
rect 42720 38010 42748 39442
rect 43456 39438 43484 39510
rect 43444 39432 43496 39438
rect 43444 39374 43496 39380
rect 43260 38956 43312 38962
rect 43260 38898 43312 38904
rect 42708 38004 42760 38010
rect 42708 37946 42760 37952
rect 42800 37868 42852 37874
rect 42800 37810 42852 37816
rect 42708 37800 42760 37806
rect 42708 37742 42760 37748
rect 42720 37466 42748 37742
rect 42708 37460 42760 37466
rect 42708 37402 42760 37408
rect 42812 37262 42840 37810
rect 43272 37806 43300 38898
rect 43456 38570 43484 39374
rect 43732 38894 43760 39782
rect 43720 38888 43772 38894
rect 43720 38830 43772 38836
rect 43916 38729 43944 41239
rect 44008 40118 44036 41386
rect 44088 41200 44140 41206
rect 44088 41142 44140 41148
rect 43996 40112 44048 40118
rect 43996 40054 44048 40060
rect 44100 39642 44128 41142
rect 44284 41070 44312 41386
rect 44272 41064 44324 41070
rect 44272 41006 44324 41012
rect 44088 39636 44140 39642
rect 44088 39578 44140 39584
rect 44376 38962 44404 44338
rect 45928 44328 45980 44334
rect 45928 44270 45980 44276
rect 44732 44260 44784 44266
rect 44732 44202 44784 44208
rect 44744 43994 44772 44202
rect 45376 44192 45428 44198
rect 45376 44134 45428 44140
rect 44732 43988 44784 43994
rect 44732 43930 44784 43936
rect 44916 43784 44968 43790
rect 44916 43726 44968 43732
rect 44456 43716 44508 43722
rect 44456 43658 44508 43664
rect 44468 42158 44496 43658
rect 44824 43240 44876 43246
rect 44824 43182 44876 43188
rect 44456 42152 44508 42158
rect 44456 42094 44508 42100
rect 44732 41676 44784 41682
rect 44732 41618 44784 41624
rect 44744 41206 44772 41618
rect 44732 41200 44784 41206
rect 44732 41142 44784 41148
rect 44836 40526 44864 43182
rect 44928 42702 44956 43726
rect 45388 43314 45416 44134
rect 45940 43314 45968 44270
rect 46020 44192 46072 44198
rect 46020 44134 46072 44140
rect 45376 43308 45428 43314
rect 45376 43250 45428 43256
rect 45928 43308 45980 43314
rect 45928 43250 45980 43256
rect 44916 42696 44968 42702
rect 44916 42638 44968 42644
rect 45284 42696 45336 42702
rect 45284 42638 45336 42644
rect 44928 42106 44956 42638
rect 45296 42362 45324 42638
rect 45284 42356 45336 42362
rect 45284 42298 45336 42304
rect 45940 42294 45968 43250
rect 46032 42906 46060 44134
rect 46020 42900 46072 42906
rect 46020 42842 46072 42848
rect 45928 42288 45980 42294
rect 45928 42230 45980 42236
rect 45836 42220 45888 42226
rect 45836 42162 45888 42168
rect 45100 42152 45152 42158
rect 44928 42100 45100 42106
rect 44928 42094 45152 42100
rect 44928 42078 45140 42094
rect 44824 40520 44876 40526
rect 44824 40462 44876 40468
rect 44824 40044 44876 40050
rect 44928 40032 44956 42078
rect 45848 42022 45876 42162
rect 45836 42016 45888 42022
rect 45836 41958 45888 41964
rect 45008 41812 45060 41818
rect 45008 41754 45060 41760
rect 45020 41138 45048 41754
rect 45940 41750 45968 42230
rect 46020 42016 46072 42022
rect 46020 41958 46072 41964
rect 46032 41818 46060 41958
rect 46020 41812 46072 41818
rect 46020 41754 46072 41760
rect 45928 41744 45980 41750
rect 45928 41686 45980 41692
rect 45836 41608 45888 41614
rect 45836 41550 45888 41556
rect 45744 41540 45796 41546
rect 45744 41482 45796 41488
rect 45756 41138 45784 41482
rect 45008 41132 45060 41138
rect 45008 41074 45060 41080
rect 45744 41132 45796 41138
rect 45744 41074 45796 41080
rect 45848 40934 45876 41550
rect 45928 41540 45980 41546
rect 45928 41482 45980 41488
rect 45100 40928 45152 40934
rect 45100 40870 45152 40876
rect 45744 40928 45796 40934
rect 45744 40870 45796 40876
rect 45836 40928 45888 40934
rect 45836 40870 45888 40876
rect 45112 40662 45140 40870
rect 45100 40656 45152 40662
rect 45100 40598 45152 40604
rect 45756 40186 45784 40870
rect 45848 40390 45876 40870
rect 45836 40384 45888 40390
rect 45836 40326 45888 40332
rect 45744 40180 45796 40186
rect 45744 40122 45796 40128
rect 44876 40004 44956 40032
rect 44824 39986 44876 39992
rect 44730 39808 44786 39817
rect 44730 39743 44786 39752
rect 44364 38956 44416 38962
rect 44364 38898 44416 38904
rect 44088 38752 44140 38758
rect 43902 38720 43958 38729
rect 44088 38694 44140 38700
rect 43902 38655 43958 38664
rect 43364 38542 43484 38570
rect 43364 37874 43392 38542
rect 44100 38486 44128 38694
rect 43444 38480 43496 38486
rect 43444 38422 43496 38428
rect 44088 38480 44140 38486
rect 44088 38422 44140 38428
rect 43456 38010 43484 38422
rect 43720 38344 43772 38350
rect 43720 38286 43772 38292
rect 43732 38214 43760 38286
rect 44744 38214 44772 39743
rect 44836 38554 44864 39986
rect 45744 39568 45796 39574
rect 45744 39510 45796 39516
rect 45284 39500 45336 39506
rect 45284 39442 45336 39448
rect 45100 39432 45152 39438
rect 45098 39400 45100 39409
rect 45152 39400 45154 39409
rect 45098 39335 45154 39344
rect 45296 39098 45324 39442
rect 45560 39432 45612 39438
rect 45560 39374 45612 39380
rect 45284 39092 45336 39098
rect 45284 39034 45336 39040
rect 44916 38752 44968 38758
rect 44916 38694 44968 38700
rect 44824 38548 44876 38554
rect 44824 38490 44876 38496
rect 43720 38208 43772 38214
rect 43720 38150 43772 38156
rect 44732 38208 44784 38214
rect 44732 38150 44784 38156
rect 44546 38040 44602 38049
rect 43444 38004 43496 38010
rect 44546 37975 44548 37984
rect 43444 37946 43496 37952
rect 44600 37975 44602 37984
rect 44548 37946 44600 37952
rect 43352 37868 43404 37874
rect 43352 37810 43404 37816
rect 43260 37800 43312 37806
rect 43260 37742 43312 37748
rect 43364 37330 43392 37810
rect 44088 37392 44140 37398
rect 44088 37334 44140 37340
rect 43352 37324 43404 37330
rect 43352 37266 43404 37272
rect 42800 37256 42852 37262
rect 42800 37198 42852 37204
rect 42248 36916 42300 36922
rect 42248 36858 42300 36864
rect 44100 36854 44128 37334
rect 44560 37312 44588 37946
rect 44928 37466 44956 38694
rect 45098 38584 45154 38593
rect 45098 38519 45154 38528
rect 45112 38282 45140 38519
rect 45284 38344 45336 38350
rect 45284 38286 45336 38292
rect 45100 38276 45152 38282
rect 45100 38218 45152 38224
rect 45296 37874 45324 38286
rect 45284 37868 45336 37874
rect 45284 37810 45336 37816
rect 45296 37738 45324 37810
rect 45284 37732 45336 37738
rect 45284 37674 45336 37680
rect 44916 37460 44968 37466
rect 44916 37402 44968 37408
rect 45572 37398 45600 39374
rect 45652 38820 45704 38826
rect 45652 38762 45704 38768
rect 45664 38554 45692 38762
rect 45652 38548 45704 38554
rect 45652 38490 45704 38496
rect 45652 38344 45704 38350
rect 45652 38286 45704 38292
rect 45664 37466 45692 38286
rect 45652 37460 45704 37466
rect 45652 37402 45704 37408
rect 45100 37392 45152 37398
rect 45020 37340 45100 37346
rect 45020 37334 45152 37340
rect 45560 37392 45612 37398
rect 45560 37334 45612 37340
rect 44640 37324 44692 37330
rect 44560 37284 44640 37312
rect 44640 37266 44692 37272
rect 44824 37324 44876 37330
rect 45020 37318 45140 37334
rect 45020 37312 45048 37318
rect 44876 37284 45048 37312
rect 44824 37266 44876 37272
rect 45756 37262 45784 39510
rect 45848 39506 45876 40326
rect 45836 39500 45888 39506
rect 45836 39442 45888 39448
rect 45940 39370 45968 41482
rect 46124 41414 46152 44338
rect 47412 44266 47440 44406
rect 52736 44328 52788 44334
rect 52736 44270 52788 44276
rect 47400 44260 47452 44266
rect 47400 44202 47452 44208
rect 48044 44260 48096 44266
rect 48044 44202 48096 44208
rect 46664 44192 46716 44198
rect 46664 44134 46716 44140
rect 46676 43926 46704 44134
rect 46664 43920 46716 43926
rect 46664 43862 46716 43868
rect 46676 43178 46704 43862
rect 47400 43784 47452 43790
rect 47400 43726 47452 43732
rect 47492 43784 47544 43790
rect 47492 43726 47544 43732
rect 47952 43784 48004 43790
rect 47952 43726 48004 43732
rect 47308 43648 47360 43654
rect 47308 43590 47360 43596
rect 47320 43314 47348 43590
rect 46848 43308 46900 43314
rect 46848 43250 46900 43256
rect 47308 43308 47360 43314
rect 47308 43250 47360 43256
rect 46664 43172 46716 43178
rect 46664 43114 46716 43120
rect 46676 42838 46704 43114
rect 46756 42900 46808 42906
rect 46756 42842 46808 42848
rect 46664 42832 46716 42838
rect 46664 42774 46716 42780
rect 46296 42628 46348 42634
rect 46296 42570 46348 42576
rect 46308 42090 46336 42570
rect 46296 42084 46348 42090
rect 46296 42026 46348 42032
rect 46676 41414 46704 42774
rect 46768 42566 46796 42842
rect 46860 42838 46888 43250
rect 46940 43240 46992 43246
rect 46940 43182 46992 43188
rect 46848 42832 46900 42838
rect 46848 42774 46900 42780
rect 46848 42696 46900 42702
rect 46848 42638 46900 42644
rect 46756 42560 46808 42566
rect 46756 42502 46808 42508
rect 46756 42220 46808 42226
rect 46756 42162 46808 42168
rect 46768 41750 46796 42162
rect 46756 41744 46808 41750
rect 46756 41686 46808 41692
rect 46032 41386 46152 41414
rect 46492 41386 46704 41414
rect 46032 41138 46060 41386
rect 46020 41132 46072 41138
rect 46020 41074 46072 41080
rect 46296 41132 46348 41138
rect 46296 41074 46348 41080
rect 46020 40996 46072 41002
rect 46020 40938 46072 40944
rect 46032 39574 46060 40938
rect 46112 40044 46164 40050
rect 46112 39986 46164 39992
rect 46124 39642 46152 39986
rect 46112 39636 46164 39642
rect 46112 39578 46164 39584
rect 46020 39568 46072 39574
rect 46020 39510 46072 39516
rect 45928 39364 45980 39370
rect 45928 39306 45980 39312
rect 46032 39098 46060 39510
rect 46308 39506 46336 41074
rect 46492 40662 46520 41386
rect 46480 40656 46532 40662
rect 46480 40598 46532 40604
rect 46492 39914 46520 40598
rect 46480 39908 46532 39914
rect 46480 39850 46532 39856
rect 46296 39500 46348 39506
rect 46296 39442 46348 39448
rect 46020 39092 46072 39098
rect 46020 39034 46072 39040
rect 46492 38894 46520 39850
rect 46664 39840 46716 39846
rect 46664 39782 46716 39788
rect 46676 39642 46704 39782
rect 46664 39636 46716 39642
rect 46664 39578 46716 39584
rect 46768 39438 46796 41686
rect 46860 41614 46888 42638
rect 46848 41608 46900 41614
rect 46848 41550 46900 41556
rect 46952 41546 46980 43182
rect 47412 42906 47440 43726
rect 47504 43450 47532 43726
rect 47492 43444 47544 43450
rect 47492 43386 47544 43392
rect 47400 42900 47452 42906
rect 47400 42842 47452 42848
rect 47504 42786 47532 43386
rect 47412 42770 47532 42786
rect 47400 42764 47532 42770
rect 47452 42758 47532 42764
rect 47400 42706 47452 42712
rect 47412 42673 47440 42706
rect 47398 42664 47454 42673
rect 47398 42599 47454 42608
rect 47412 41818 47440 42599
rect 47768 42220 47820 42226
rect 47768 42162 47820 42168
rect 47400 41812 47452 41818
rect 47400 41754 47452 41760
rect 47584 41608 47636 41614
rect 47584 41550 47636 41556
rect 46940 41540 46992 41546
rect 46940 41482 46992 41488
rect 46952 41070 46980 41482
rect 46940 41064 46992 41070
rect 46940 41006 46992 41012
rect 47216 40996 47268 41002
rect 47216 40938 47268 40944
rect 47228 40458 47256 40938
rect 47596 40458 47624 41550
rect 47780 40662 47808 42162
rect 47860 41676 47912 41682
rect 47860 41618 47912 41624
rect 47768 40656 47820 40662
rect 47872 40633 47900 41618
rect 47964 40662 47992 43726
rect 48056 42090 48084 44202
rect 50918 44092 51226 44101
rect 50918 44090 50924 44092
rect 50980 44090 51004 44092
rect 51060 44090 51084 44092
rect 51140 44090 51164 44092
rect 51220 44090 51226 44092
rect 50980 44038 50982 44090
rect 51162 44038 51164 44090
rect 50918 44036 50924 44038
rect 50980 44036 51004 44038
rect 51060 44036 51084 44038
rect 51140 44036 51164 44038
rect 51220 44036 51226 44038
rect 50918 44027 51226 44036
rect 52748 43858 52776 44270
rect 53840 44192 53892 44198
rect 53840 44134 53892 44140
rect 52552 43852 52604 43858
rect 52552 43794 52604 43800
rect 52736 43852 52788 43858
rect 52736 43794 52788 43800
rect 48228 43648 48280 43654
rect 48228 43590 48280 43596
rect 51908 43648 51960 43654
rect 51908 43590 51960 43596
rect 48240 42906 48268 43590
rect 49998 43548 50306 43557
rect 49998 43546 50004 43548
rect 50060 43546 50084 43548
rect 50140 43546 50164 43548
rect 50220 43546 50244 43548
rect 50300 43546 50306 43548
rect 50060 43494 50062 43546
rect 50242 43494 50244 43546
rect 49998 43492 50004 43494
rect 50060 43492 50084 43494
rect 50140 43492 50164 43494
rect 50220 43492 50244 43494
rect 50300 43492 50306 43494
rect 49998 43483 50306 43492
rect 49516 43444 49568 43450
rect 49516 43386 49568 43392
rect 48964 43172 49016 43178
rect 48964 43114 49016 43120
rect 48228 42900 48280 42906
rect 48228 42842 48280 42848
rect 48412 42696 48464 42702
rect 48412 42638 48464 42644
rect 48044 42084 48096 42090
rect 48044 42026 48096 42032
rect 48320 42084 48372 42090
rect 48320 42026 48372 42032
rect 48136 42016 48188 42022
rect 48136 41958 48188 41964
rect 48148 41818 48176 41958
rect 48136 41812 48188 41818
rect 48136 41754 48188 41760
rect 48136 41540 48188 41546
rect 48136 41482 48188 41488
rect 47952 40656 48004 40662
rect 47768 40598 47820 40604
rect 47858 40624 47914 40633
rect 47952 40598 48004 40604
rect 47858 40559 47860 40568
rect 47912 40559 47914 40568
rect 47860 40530 47912 40536
rect 47216 40452 47268 40458
rect 47216 40394 47268 40400
rect 47584 40452 47636 40458
rect 47584 40394 47636 40400
rect 46756 39432 46808 39438
rect 46756 39374 46808 39380
rect 48148 39370 48176 41482
rect 48332 41070 48360 42026
rect 48424 41614 48452 42638
rect 48504 42016 48556 42022
rect 48504 41958 48556 41964
rect 48516 41818 48544 41958
rect 48504 41812 48556 41818
rect 48504 41754 48556 41760
rect 48412 41608 48464 41614
rect 48412 41550 48464 41556
rect 48504 41200 48556 41206
rect 48504 41142 48556 41148
rect 48320 41064 48372 41070
rect 48320 41006 48372 41012
rect 48228 40928 48280 40934
rect 48228 40870 48280 40876
rect 48240 40633 48268 40870
rect 48226 40624 48282 40633
rect 48226 40559 48282 40568
rect 48332 39574 48360 41006
rect 48516 40390 48544 41142
rect 48976 40934 49004 43114
rect 49148 42220 49200 42226
rect 49148 42162 49200 42168
rect 49160 41614 49188 42162
rect 49148 41608 49200 41614
rect 49148 41550 49200 41556
rect 48688 40928 48740 40934
rect 48688 40870 48740 40876
rect 48964 40928 49016 40934
rect 48964 40870 49016 40876
rect 48504 40384 48556 40390
rect 48504 40326 48556 40332
rect 48596 40384 48648 40390
rect 48596 40326 48648 40332
rect 48412 39636 48464 39642
rect 48412 39578 48464 39584
rect 48320 39568 48372 39574
rect 48320 39510 48372 39516
rect 48424 39438 48452 39578
rect 48516 39522 48544 40326
rect 48608 40186 48636 40326
rect 48596 40180 48648 40186
rect 48596 40122 48648 40128
rect 48516 39494 48636 39522
rect 48412 39432 48464 39438
rect 48412 39374 48464 39380
rect 48136 39364 48188 39370
rect 48136 39306 48188 39312
rect 47400 39296 47452 39302
rect 47400 39238 47452 39244
rect 47124 38956 47176 38962
rect 47124 38898 47176 38904
rect 46480 38888 46532 38894
rect 46480 38830 46532 38836
rect 46940 38752 46992 38758
rect 46940 38694 46992 38700
rect 46952 37806 46980 38694
rect 47136 38350 47164 38898
rect 47412 38554 47440 39238
rect 48148 38894 48176 39306
rect 48424 38894 48452 39374
rect 47860 38888 47912 38894
rect 47860 38830 47912 38836
rect 48136 38888 48188 38894
rect 48136 38830 48188 38836
rect 48412 38888 48464 38894
rect 48412 38830 48464 38836
rect 47584 38820 47636 38826
rect 47584 38762 47636 38768
rect 47596 38554 47624 38762
rect 47872 38758 47900 38830
rect 47860 38752 47912 38758
rect 47860 38694 47912 38700
rect 47400 38548 47452 38554
rect 47400 38490 47452 38496
rect 47584 38548 47636 38554
rect 47584 38490 47636 38496
rect 47872 38486 47900 38694
rect 48318 38584 48374 38593
rect 48318 38519 48374 38528
rect 47860 38480 47912 38486
rect 47860 38422 47912 38428
rect 47124 38344 47176 38350
rect 47124 38286 47176 38292
rect 47768 38344 47820 38350
rect 47768 38286 47820 38292
rect 46940 37800 46992 37806
rect 46940 37742 46992 37748
rect 46020 37732 46072 37738
rect 46020 37674 46072 37680
rect 46032 37466 46060 37674
rect 46940 37664 46992 37670
rect 46940 37606 46992 37612
rect 46020 37460 46072 37466
rect 46020 37402 46072 37408
rect 46952 37398 46980 37606
rect 46940 37392 46992 37398
rect 46940 37334 46992 37340
rect 45744 37256 45796 37262
rect 45744 37198 45796 37204
rect 46756 37188 46808 37194
rect 46756 37130 46808 37136
rect 44088 36848 44140 36854
rect 44088 36790 44140 36796
rect 46768 36786 46796 37130
rect 47136 37126 47164 38286
rect 47780 37466 47808 38286
rect 48332 37874 48360 38519
rect 48608 38350 48636 39494
rect 48700 38962 48728 40870
rect 48976 39914 49004 40870
rect 49160 40526 49188 41550
rect 49528 41206 49556 43386
rect 51264 43308 51316 43314
rect 51264 43250 51316 43256
rect 50918 43004 51226 43013
rect 50918 43002 50924 43004
rect 50980 43002 51004 43004
rect 51060 43002 51084 43004
rect 51140 43002 51164 43004
rect 51220 43002 51226 43004
rect 50980 42950 50982 43002
rect 51162 42950 51164 43002
rect 50918 42948 50924 42950
rect 50980 42948 51004 42950
rect 51060 42948 51084 42950
rect 51140 42948 51164 42950
rect 51220 42948 51226 42950
rect 50918 42939 51226 42948
rect 49998 42460 50306 42469
rect 49998 42458 50004 42460
rect 50060 42458 50084 42460
rect 50140 42458 50164 42460
rect 50220 42458 50244 42460
rect 50300 42458 50306 42460
rect 50060 42406 50062 42458
rect 50242 42406 50244 42458
rect 49998 42404 50004 42406
rect 50060 42404 50084 42406
rect 50140 42404 50164 42406
rect 50220 42404 50244 42406
rect 50300 42404 50306 42406
rect 49998 42395 50306 42404
rect 49700 42356 49752 42362
rect 49700 42298 49752 42304
rect 49516 41200 49568 41206
rect 49516 41142 49568 41148
rect 49608 41064 49660 41070
rect 49608 41006 49660 41012
rect 49056 40520 49108 40526
rect 49056 40462 49108 40468
rect 49148 40520 49200 40526
rect 49148 40462 49200 40468
rect 48964 39908 49016 39914
rect 48964 39850 49016 39856
rect 48872 39568 48924 39574
rect 48872 39510 48924 39516
rect 48780 39500 48832 39506
rect 48780 39442 48832 39448
rect 48688 38956 48740 38962
rect 48688 38898 48740 38904
rect 48792 38554 48820 39442
rect 48884 38593 48912 39510
rect 49068 39098 49096 40462
rect 49240 40452 49292 40458
rect 49240 40394 49292 40400
rect 49056 39092 49108 39098
rect 49056 39034 49108 39040
rect 49252 38962 49280 40394
rect 49620 40186 49648 41006
rect 49712 40662 49740 42298
rect 49884 42084 49936 42090
rect 49884 42026 49936 42032
rect 49792 42016 49844 42022
rect 49792 41958 49844 41964
rect 49804 41002 49832 41958
rect 49792 40996 49844 41002
rect 49792 40938 49844 40944
rect 49700 40656 49752 40662
rect 49700 40598 49752 40604
rect 49608 40180 49660 40186
rect 49608 40122 49660 40128
rect 49712 40050 49740 40598
rect 49792 40588 49844 40594
rect 49792 40530 49844 40536
rect 49804 40497 49832 40530
rect 49790 40488 49846 40497
rect 49896 40458 49924 42026
rect 50436 42016 50488 42022
rect 50436 41958 50488 41964
rect 50712 42016 50764 42022
rect 50712 41958 50764 41964
rect 50448 41818 50476 41958
rect 50436 41812 50488 41818
rect 50436 41754 50488 41760
rect 50344 41744 50396 41750
rect 50344 41686 50396 41692
rect 49998 41372 50306 41381
rect 49998 41370 50004 41372
rect 50060 41370 50084 41372
rect 50140 41370 50164 41372
rect 50220 41370 50244 41372
rect 50300 41370 50306 41372
rect 50060 41318 50062 41370
rect 50242 41318 50244 41370
rect 49998 41316 50004 41318
rect 50060 41316 50084 41318
rect 50140 41316 50164 41318
rect 50220 41316 50244 41318
rect 50300 41316 50306 41318
rect 49998 41307 50306 41316
rect 50356 41002 50384 41686
rect 50724 41614 50752 41958
rect 50918 41916 51226 41925
rect 50918 41914 50924 41916
rect 50980 41914 51004 41916
rect 51060 41914 51084 41916
rect 51140 41914 51164 41916
rect 51220 41914 51226 41916
rect 50980 41862 50982 41914
rect 51162 41862 51164 41914
rect 50918 41860 50924 41862
rect 50980 41860 51004 41862
rect 51060 41860 51084 41862
rect 51140 41860 51164 41862
rect 51220 41860 51226 41862
rect 50918 41851 51226 41860
rect 50712 41608 50764 41614
rect 50712 41550 50764 41556
rect 50344 40996 50396 41002
rect 50344 40938 50396 40944
rect 50724 40594 50752 41550
rect 50896 41132 50948 41138
rect 50896 41074 50948 41080
rect 50908 41041 50936 41074
rect 50894 41032 50950 41041
rect 50894 40967 50950 40976
rect 50918 40828 51226 40837
rect 50918 40826 50924 40828
rect 50980 40826 51004 40828
rect 51060 40826 51084 40828
rect 51140 40826 51164 40828
rect 51220 40826 51226 40828
rect 50980 40774 50982 40826
rect 51162 40774 51164 40826
rect 50918 40772 50924 40774
rect 50980 40772 51004 40774
rect 51060 40772 51084 40774
rect 51140 40772 51164 40774
rect 51220 40772 51226 40774
rect 50918 40763 51226 40772
rect 50712 40588 50764 40594
rect 50712 40530 50764 40536
rect 50436 40520 50488 40526
rect 50436 40462 50488 40468
rect 49790 40423 49846 40432
rect 49884 40452 49936 40458
rect 49884 40394 49936 40400
rect 49998 40284 50306 40293
rect 49998 40282 50004 40284
rect 50060 40282 50084 40284
rect 50140 40282 50164 40284
rect 50220 40282 50244 40284
rect 50300 40282 50306 40284
rect 50060 40230 50062 40282
rect 50242 40230 50244 40282
rect 49998 40228 50004 40230
rect 50060 40228 50084 40230
rect 50140 40228 50164 40230
rect 50220 40228 50244 40230
rect 50300 40228 50306 40230
rect 49998 40219 50306 40228
rect 50448 40118 50476 40462
rect 50620 40384 50672 40390
rect 50620 40326 50672 40332
rect 49884 40112 49936 40118
rect 49884 40054 49936 40060
rect 50436 40112 50488 40118
rect 50436 40054 50488 40060
rect 49700 40044 49752 40050
rect 49700 39986 49752 39992
rect 49896 39846 49924 40054
rect 49884 39840 49936 39846
rect 49884 39782 49936 39788
rect 49976 39840 50028 39846
rect 49976 39782 50028 39788
rect 50252 39840 50304 39846
rect 50252 39782 50304 39788
rect 49896 39642 49924 39782
rect 49988 39642 50016 39782
rect 49884 39636 49936 39642
rect 49884 39578 49936 39584
rect 49976 39636 50028 39642
rect 49976 39578 50028 39584
rect 50264 39574 50292 39782
rect 50632 39574 50660 40326
rect 51276 40202 51304 43250
rect 51540 43104 51592 43110
rect 51540 43046 51592 43052
rect 51552 42906 51580 43046
rect 51540 42900 51592 42906
rect 51540 42842 51592 42848
rect 51920 42702 51948 43590
rect 52564 43450 52592 43794
rect 52552 43444 52604 43450
rect 52552 43386 52604 43392
rect 52552 43308 52604 43314
rect 52552 43250 52604 43256
rect 52460 43104 52512 43110
rect 52460 43046 52512 43052
rect 52472 42906 52500 43046
rect 52460 42900 52512 42906
rect 52460 42842 52512 42848
rect 51724 42696 51776 42702
rect 51724 42638 51776 42644
rect 51908 42696 51960 42702
rect 51908 42638 51960 42644
rect 52460 42696 52512 42702
rect 52460 42638 52512 42644
rect 51540 42628 51592 42634
rect 51540 42570 51592 42576
rect 51356 42084 51408 42090
rect 51356 42026 51408 42032
rect 51368 41546 51396 42026
rect 51356 41540 51408 41546
rect 51356 41482 51408 41488
rect 51368 41274 51396 41482
rect 51356 41268 51408 41274
rect 51356 41210 51408 41216
rect 51552 40458 51580 42570
rect 51736 42362 51764 42638
rect 51920 42566 51948 42638
rect 51908 42560 51960 42566
rect 51908 42502 51960 42508
rect 52472 42362 52500 42638
rect 51632 42356 51684 42362
rect 51632 42298 51684 42304
rect 51724 42356 51776 42362
rect 51724 42298 51776 42304
rect 52460 42356 52512 42362
rect 52460 42298 52512 42304
rect 51644 42242 51672 42298
rect 51644 42226 51764 42242
rect 51644 42220 51776 42226
rect 51644 42214 51724 42220
rect 51724 42162 51776 42168
rect 52564 42158 52592 43250
rect 52644 42220 52696 42226
rect 52644 42162 52696 42168
rect 52368 42152 52420 42158
rect 52368 42094 52420 42100
rect 52552 42152 52604 42158
rect 52552 42094 52604 42100
rect 52380 41818 52408 42094
rect 52656 42022 52684 42162
rect 52460 42016 52512 42022
rect 52644 42016 52696 42022
rect 52512 41976 52592 42004
rect 52460 41958 52512 41964
rect 52368 41812 52420 41818
rect 52368 41754 52420 41760
rect 52368 41608 52420 41614
rect 52368 41550 52420 41556
rect 52184 40996 52236 41002
rect 52184 40938 52236 40944
rect 52196 40594 52224 40938
rect 52184 40588 52236 40594
rect 52184 40530 52236 40536
rect 51540 40452 51592 40458
rect 51540 40394 51592 40400
rect 51276 40186 51396 40202
rect 51276 40180 51408 40186
rect 51276 40174 51356 40180
rect 51356 40122 51408 40128
rect 50712 39908 50764 39914
rect 50712 39850 50764 39856
rect 50252 39568 50304 39574
rect 50252 39510 50304 39516
rect 50620 39568 50672 39574
rect 50620 39510 50672 39516
rect 50724 39438 50752 39850
rect 50918 39740 51226 39749
rect 50918 39738 50924 39740
rect 50980 39738 51004 39740
rect 51060 39738 51084 39740
rect 51140 39738 51164 39740
rect 51220 39738 51226 39740
rect 50980 39686 50982 39738
rect 51162 39686 51164 39738
rect 50918 39684 50924 39686
rect 50980 39684 51004 39686
rect 51060 39684 51084 39686
rect 51140 39684 51164 39686
rect 51220 39684 51226 39686
rect 50918 39675 51226 39684
rect 51368 39574 51396 40122
rect 51552 40118 51580 40394
rect 51540 40112 51592 40118
rect 51540 40054 51592 40060
rect 52092 39908 52144 39914
rect 52092 39850 52144 39856
rect 51356 39568 51408 39574
rect 51356 39510 51408 39516
rect 50712 39432 50764 39438
rect 50712 39374 50764 39380
rect 50804 39364 50856 39370
rect 50804 39306 50856 39312
rect 49998 39196 50306 39205
rect 49998 39194 50004 39196
rect 50060 39194 50084 39196
rect 50140 39194 50164 39196
rect 50220 39194 50244 39196
rect 50300 39194 50306 39196
rect 50060 39142 50062 39194
rect 50242 39142 50244 39194
rect 49998 39140 50004 39142
rect 50060 39140 50084 39142
rect 50140 39140 50164 39142
rect 50220 39140 50244 39142
rect 50300 39140 50306 39142
rect 49998 39131 50306 39140
rect 49240 38956 49292 38962
rect 49240 38898 49292 38904
rect 49884 38752 49936 38758
rect 49884 38694 49936 38700
rect 50344 38752 50396 38758
rect 50344 38694 50396 38700
rect 48870 38584 48926 38593
rect 48688 38548 48740 38554
rect 48688 38490 48740 38496
rect 48780 38548 48832 38554
rect 48870 38519 48926 38528
rect 48780 38490 48832 38496
rect 48596 38344 48648 38350
rect 48596 38286 48648 38292
rect 48320 37868 48372 37874
rect 48320 37810 48372 37816
rect 48412 37868 48464 37874
rect 48464 37828 48544 37856
rect 48412 37810 48464 37816
rect 48320 37732 48372 37738
rect 48372 37692 48452 37720
rect 48320 37674 48372 37680
rect 48228 37664 48280 37670
rect 48228 37606 48280 37612
rect 48240 37466 48268 37606
rect 47768 37460 47820 37466
rect 47768 37402 47820 37408
rect 48228 37460 48280 37466
rect 48228 37402 48280 37408
rect 48424 37369 48452 37692
rect 48516 37466 48544 37828
rect 48504 37460 48556 37466
rect 48504 37402 48556 37408
rect 48410 37360 48466 37369
rect 48410 37295 48466 37304
rect 48608 37262 48636 38286
rect 47216 37256 47268 37262
rect 47216 37198 47268 37204
rect 48596 37256 48648 37262
rect 48596 37198 48648 37204
rect 47124 37120 47176 37126
rect 47124 37062 47176 37068
rect 47228 36922 47256 37198
rect 48608 36922 48636 37198
rect 48700 37194 48728 38490
rect 49896 38486 49924 38694
rect 49974 38584 50030 38593
rect 49974 38519 50030 38528
rect 49988 38486 50016 38519
rect 49884 38480 49936 38486
rect 49884 38422 49936 38428
rect 49976 38480 50028 38486
rect 49976 38422 50028 38428
rect 49998 38108 50306 38117
rect 49998 38106 50004 38108
rect 50060 38106 50084 38108
rect 50140 38106 50164 38108
rect 50220 38106 50244 38108
rect 50300 38106 50306 38108
rect 50060 38054 50062 38106
rect 50242 38054 50244 38106
rect 49998 38052 50004 38054
rect 50060 38052 50084 38054
rect 50140 38052 50164 38054
rect 50220 38052 50244 38054
rect 50300 38052 50306 38054
rect 49998 38043 50306 38052
rect 50356 37856 50384 38694
rect 50816 38010 50844 39306
rect 50918 38652 51226 38661
rect 50918 38650 50924 38652
rect 50980 38650 51004 38652
rect 51060 38650 51084 38652
rect 51140 38650 51164 38652
rect 51220 38650 51226 38652
rect 50980 38598 50982 38650
rect 51162 38598 51164 38650
rect 50918 38596 50924 38598
rect 50980 38596 51004 38598
rect 51060 38596 51084 38598
rect 51140 38596 51164 38598
rect 51220 38596 51226 38598
rect 50918 38587 51226 38596
rect 51172 38480 51224 38486
rect 51092 38440 51172 38468
rect 51092 38350 51120 38440
rect 51172 38422 51224 38428
rect 51080 38344 51132 38350
rect 51080 38286 51132 38292
rect 51264 38276 51316 38282
rect 51264 38218 51316 38224
rect 50804 38004 50856 38010
rect 50804 37946 50856 37952
rect 50264 37828 50384 37856
rect 49332 37800 49384 37806
rect 49332 37742 49384 37748
rect 49344 37398 49372 37742
rect 50264 37466 50292 37828
rect 50344 37732 50396 37738
rect 50344 37674 50396 37680
rect 50356 37466 50384 37674
rect 50918 37564 51226 37573
rect 50918 37562 50924 37564
rect 50980 37562 51004 37564
rect 51060 37562 51084 37564
rect 51140 37562 51164 37564
rect 51220 37562 51226 37564
rect 50980 37510 50982 37562
rect 51162 37510 51164 37562
rect 50918 37508 50924 37510
rect 50980 37508 51004 37510
rect 51060 37508 51084 37510
rect 51140 37508 51164 37510
rect 51220 37508 51226 37510
rect 50918 37499 51226 37508
rect 51276 37466 51304 38218
rect 51368 37874 51396 39510
rect 52104 39506 52132 39850
rect 52196 39574 52224 40530
rect 52380 39642 52408 41550
rect 52564 41478 52592 41976
rect 52644 41958 52696 41964
rect 52460 41472 52512 41478
rect 52460 41414 52512 41420
rect 52552 41472 52604 41478
rect 52552 41414 52604 41420
rect 52472 40662 52500 41414
rect 52460 40656 52512 40662
rect 52460 40598 52512 40604
rect 52368 39636 52420 39642
rect 52368 39578 52420 39584
rect 52184 39568 52236 39574
rect 52564 39545 52592 41414
rect 52656 41138 52684 41958
rect 52644 41132 52696 41138
rect 52644 41074 52696 41080
rect 52644 40384 52696 40390
rect 52644 40326 52696 40332
rect 52184 39510 52236 39516
rect 52550 39536 52606 39545
rect 52092 39500 52144 39506
rect 52656 39506 52684 40326
rect 52748 39828 52776 43794
rect 53196 43648 53248 43654
rect 53196 43590 53248 43596
rect 53208 43178 53236 43590
rect 53852 43246 53880 44134
rect 66352 43852 66404 43858
rect 66352 43794 66404 43800
rect 53840 43240 53892 43246
rect 53840 43182 53892 43188
rect 53196 43172 53248 43178
rect 53196 43114 53248 43120
rect 52828 42696 52880 42702
rect 52828 42638 52880 42644
rect 52840 41478 52868 42638
rect 52920 42560 52972 42566
rect 52920 42502 52972 42508
rect 52932 41614 52960 42502
rect 53208 42362 53236 43114
rect 53380 43104 53432 43110
rect 53380 43046 53432 43052
rect 53196 42356 53248 42362
rect 53196 42298 53248 42304
rect 53208 42090 53236 42298
rect 53392 42294 53420 43046
rect 53380 42288 53432 42294
rect 53380 42230 53432 42236
rect 53392 42158 53420 42230
rect 53852 42158 53880 43182
rect 60648 43104 60700 43110
rect 60648 43046 60700 43052
rect 54024 42832 54076 42838
rect 54024 42774 54076 42780
rect 53932 42220 53984 42226
rect 53932 42162 53984 42168
rect 53380 42152 53432 42158
rect 53380 42094 53432 42100
rect 53840 42152 53892 42158
rect 53840 42094 53892 42100
rect 53196 42084 53248 42090
rect 53196 42026 53248 42032
rect 52920 41608 52972 41614
rect 52920 41550 52972 41556
rect 53840 41608 53892 41614
rect 53840 41550 53892 41556
rect 52932 41478 52960 41550
rect 52828 41472 52880 41478
rect 52828 41414 52880 41420
rect 52920 41472 52972 41478
rect 52920 41414 52972 41420
rect 52828 39840 52880 39846
rect 52748 39800 52828 39828
rect 52748 39642 52776 39800
rect 52828 39782 52880 39788
rect 52736 39636 52788 39642
rect 52736 39578 52788 39584
rect 52828 39568 52880 39574
rect 52826 39536 52828 39545
rect 52880 39536 52882 39545
rect 52550 39471 52606 39480
rect 52644 39500 52696 39506
rect 52092 39442 52144 39448
rect 52826 39471 52882 39480
rect 52644 39442 52696 39448
rect 51448 38888 51500 38894
rect 52104 38865 52132 39442
rect 51448 38830 51500 38836
rect 52090 38856 52146 38865
rect 51460 38554 51488 38830
rect 52090 38791 52146 38800
rect 51448 38548 51500 38554
rect 51448 38490 51500 38496
rect 51460 38214 51488 38490
rect 52932 38350 52960 41414
rect 53104 41268 53156 41274
rect 53104 41210 53156 41216
rect 53116 40662 53144 41210
rect 53472 40928 53524 40934
rect 53472 40870 53524 40876
rect 53656 40928 53708 40934
rect 53852 40882 53880 41550
rect 53944 41138 53972 42162
rect 54036 42090 54064 42774
rect 59268 42356 59320 42362
rect 59268 42298 59320 42304
rect 58070 42256 58126 42265
rect 58070 42191 58126 42200
rect 54024 42084 54076 42090
rect 54024 42026 54076 42032
rect 55772 42084 55824 42090
rect 55772 42026 55824 42032
rect 54036 41274 54064 42026
rect 55312 41608 55364 41614
rect 55312 41550 55364 41556
rect 55036 41472 55088 41478
rect 55036 41414 55088 41420
rect 54024 41268 54076 41274
rect 54024 41210 54076 41216
rect 53932 41132 53984 41138
rect 53932 41074 53984 41080
rect 53708 40876 53880 40882
rect 53656 40870 53880 40876
rect 53932 40928 53984 40934
rect 53932 40870 53984 40876
rect 53104 40656 53156 40662
rect 53104 40598 53156 40604
rect 53116 39914 53144 40598
rect 53484 40050 53512 40870
rect 53668 40854 53880 40870
rect 53852 40526 53880 40854
rect 53840 40520 53892 40526
rect 53840 40462 53892 40468
rect 53944 40390 53972 40870
rect 54036 40662 54064 41210
rect 54116 41132 54168 41138
rect 54116 41074 54168 41080
rect 54128 40934 54156 41074
rect 54760 41064 54812 41070
rect 54760 41006 54812 41012
rect 54116 40928 54168 40934
rect 54116 40870 54168 40876
rect 54668 40928 54720 40934
rect 54668 40870 54720 40876
rect 54024 40656 54076 40662
rect 54024 40598 54076 40604
rect 54576 40520 54628 40526
rect 54576 40462 54628 40468
rect 53932 40384 53984 40390
rect 53932 40326 53984 40332
rect 54588 40186 54616 40462
rect 54576 40180 54628 40186
rect 54576 40122 54628 40128
rect 54680 40050 54708 40870
rect 53472 40044 53524 40050
rect 53472 39986 53524 39992
rect 54668 40044 54720 40050
rect 54668 39986 54720 39992
rect 53104 39908 53156 39914
rect 53024 39868 53104 39896
rect 53024 38826 53052 39868
rect 53104 39850 53156 39856
rect 54484 39840 54536 39846
rect 54484 39782 54536 39788
rect 53564 39432 53616 39438
rect 53564 39374 53616 39380
rect 53196 39296 53248 39302
rect 53196 39238 53248 39244
rect 53012 38820 53064 38826
rect 53012 38762 53064 38768
rect 51816 38344 51868 38350
rect 51816 38286 51868 38292
rect 52920 38344 52972 38350
rect 52920 38286 52972 38292
rect 51448 38208 51500 38214
rect 51448 38150 51500 38156
rect 51828 38010 51856 38286
rect 52276 38208 52328 38214
rect 52276 38150 52328 38156
rect 51816 38004 51868 38010
rect 51816 37946 51868 37952
rect 51356 37868 51408 37874
rect 51356 37810 51408 37816
rect 50252 37460 50304 37466
rect 50252 37402 50304 37408
rect 50344 37460 50396 37466
rect 50344 37402 50396 37408
rect 51264 37460 51316 37466
rect 51264 37402 51316 37408
rect 51828 37398 51856 37946
rect 52288 37466 52316 38150
rect 52552 37732 52604 37738
rect 52552 37674 52604 37680
rect 52564 37482 52592 37674
rect 52564 37466 52776 37482
rect 52276 37460 52328 37466
rect 52276 37402 52328 37408
rect 52564 37460 52788 37466
rect 52564 37454 52736 37460
rect 49332 37392 49384 37398
rect 49332 37334 49384 37340
rect 51816 37392 51868 37398
rect 51816 37334 51868 37340
rect 48688 37188 48740 37194
rect 48688 37130 48740 37136
rect 49998 37020 50306 37029
rect 49998 37018 50004 37020
rect 50060 37018 50084 37020
rect 50140 37018 50164 37020
rect 50220 37018 50244 37020
rect 50300 37018 50306 37020
rect 50060 36966 50062 37018
rect 50242 36966 50244 37018
rect 49998 36964 50004 36966
rect 50060 36964 50084 36966
rect 50140 36964 50164 36966
rect 50220 36964 50244 36966
rect 50300 36964 50306 36966
rect 49998 36955 50306 36964
rect 47216 36916 47268 36922
rect 47216 36858 47268 36864
rect 48596 36916 48648 36922
rect 48596 36858 48648 36864
rect 46756 36780 46808 36786
rect 46756 36722 46808 36728
rect 41694 36680 41750 36689
rect 41694 36615 41750 36624
rect 52564 36514 52592 37454
rect 52736 37402 52788 37408
rect 52932 37330 52960 38286
rect 53024 37806 53052 38762
rect 53208 38554 53236 39238
rect 53576 38758 53604 39374
rect 53656 38820 53708 38826
rect 53656 38762 53708 38768
rect 53564 38752 53616 38758
rect 53564 38694 53616 38700
rect 53196 38548 53248 38554
rect 53196 38490 53248 38496
rect 53380 38412 53432 38418
rect 53380 38354 53432 38360
rect 53392 38214 53420 38354
rect 53380 38208 53432 38214
rect 53380 38150 53432 38156
rect 53012 37800 53064 37806
rect 53012 37742 53064 37748
rect 53576 37466 53604 38694
rect 53668 38554 53696 38762
rect 53656 38548 53708 38554
rect 53656 38490 53708 38496
rect 54496 38486 54524 39782
rect 54680 39506 54708 39986
rect 54772 39574 54800 41006
rect 55048 41002 55076 41414
rect 55036 40996 55088 41002
rect 55036 40938 55088 40944
rect 55128 40996 55180 41002
rect 55128 40938 55180 40944
rect 55140 40662 55168 40938
rect 55128 40656 55180 40662
rect 55128 40598 55180 40604
rect 55036 40384 55088 40390
rect 55036 40326 55088 40332
rect 55048 40118 55076 40326
rect 55036 40112 55088 40118
rect 55036 40054 55088 40060
rect 55140 40066 55168 40598
rect 55140 40038 55260 40066
rect 54760 39568 54812 39574
rect 54760 39510 54812 39516
rect 54668 39500 54720 39506
rect 54668 39442 54720 39448
rect 54024 38480 54076 38486
rect 53760 38418 53972 38434
rect 54024 38422 54076 38428
rect 54484 38480 54536 38486
rect 54484 38422 54536 38428
rect 53760 38412 53984 38418
rect 53760 38406 53932 38412
rect 53656 37664 53708 37670
rect 53760 37618 53788 38406
rect 53932 38354 53984 38360
rect 53840 38208 53892 38214
rect 54036 38196 54064 38422
rect 54680 38350 54708 39442
rect 55232 38758 55260 40038
rect 55324 39846 55352 41550
rect 55784 41041 55812 42026
rect 56324 42016 56376 42022
rect 56324 41958 56376 41964
rect 56336 41414 56364 41958
rect 56508 41608 56560 41614
rect 56508 41550 56560 41556
rect 56244 41386 56364 41414
rect 55770 41032 55826 41041
rect 55770 40967 55826 40976
rect 55588 40520 55640 40526
rect 55588 40462 55640 40468
rect 56048 40520 56100 40526
rect 56048 40462 56100 40468
rect 55600 40186 55628 40462
rect 55588 40180 55640 40186
rect 55588 40122 55640 40128
rect 56060 39914 56088 40462
rect 56244 40050 56272 41386
rect 56520 41274 56548 41550
rect 57428 41540 57480 41546
rect 57428 41482 57480 41488
rect 56508 41268 56560 41274
rect 56508 41210 56560 41216
rect 56232 40044 56284 40050
rect 56232 39986 56284 39992
rect 56048 39908 56100 39914
rect 56048 39850 56100 39856
rect 55312 39840 55364 39846
rect 55312 39782 55364 39788
rect 55956 39432 56008 39438
rect 55956 39374 56008 39380
rect 55312 39296 55364 39302
rect 55312 39238 55364 39244
rect 55324 38826 55352 39238
rect 55312 38820 55364 38826
rect 55312 38762 55364 38768
rect 55772 38820 55824 38826
rect 55772 38762 55824 38768
rect 55220 38752 55272 38758
rect 55220 38694 55272 38700
rect 55218 38448 55274 38457
rect 55784 38418 55812 38762
rect 55218 38383 55220 38392
rect 55272 38383 55274 38392
rect 55772 38412 55824 38418
rect 55220 38354 55272 38360
rect 55772 38354 55824 38360
rect 54668 38344 54720 38350
rect 54668 38286 54720 38292
rect 53892 38168 54064 38196
rect 53840 38150 53892 38156
rect 53708 37612 53788 37618
rect 53656 37606 53788 37612
rect 53668 37590 53788 37606
rect 53196 37460 53248 37466
rect 53196 37402 53248 37408
rect 53564 37460 53616 37466
rect 53564 37402 53616 37408
rect 52920 37324 52972 37330
rect 52920 37266 52972 37272
rect 53208 37194 53236 37402
rect 53760 37194 53788 37590
rect 53852 37369 53880 38150
rect 54680 37874 54708 38286
rect 54668 37868 54720 37874
rect 54668 37810 54720 37816
rect 54300 37732 54352 37738
rect 54300 37674 54352 37680
rect 54312 37466 54340 37674
rect 54300 37460 54352 37466
rect 54300 37402 54352 37408
rect 53838 37360 53894 37369
rect 53838 37295 53894 37304
rect 53196 37188 53248 37194
rect 53196 37130 53248 37136
rect 53748 37188 53800 37194
rect 53748 37130 53800 37136
rect 54680 37126 54708 37810
rect 55232 37806 55260 38354
rect 55968 37942 55996 39374
rect 56244 39302 56272 39986
rect 56520 39982 56548 41210
rect 57440 41070 57468 41482
rect 58084 41206 58112 42191
rect 58072 41200 58124 41206
rect 58072 41142 58124 41148
rect 56692 41064 56744 41070
rect 56598 41032 56654 41041
rect 56692 41006 56744 41012
rect 57428 41064 57480 41070
rect 57428 41006 57480 41012
rect 56598 40967 56600 40976
rect 56652 40967 56654 40976
rect 56600 40938 56652 40944
rect 56508 39976 56560 39982
rect 56508 39918 56560 39924
rect 56324 39432 56376 39438
rect 56324 39374 56376 39380
rect 56232 39296 56284 39302
rect 56232 39238 56284 39244
rect 56048 38956 56100 38962
rect 56048 38898 56100 38904
rect 55956 37936 56008 37942
rect 55956 37878 56008 37884
rect 56060 37806 56088 38898
rect 56244 37874 56272 39238
rect 56336 38962 56364 39374
rect 56324 38956 56376 38962
rect 56324 38898 56376 38904
rect 56232 37868 56284 37874
rect 56232 37810 56284 37816
rect 55220 37800 55272 37806
rect 55220 37742 55272 37748
rect 56048 37800 56100 37806
rect 56048 37742 56100 37748
rect 56060 37330 56088 37742
rect 56048 37324 56100 37330
rect 56048 37266 56100 37272
rect 54668 37120 54720 37126
rect 54668 37062 54720 37068
rect 52552 36508 52604 36514
rect 52552 36450 52604 36456
rect 42706 36408 42762 36417
rect 42706 36343 42762 36352
rect 40130 35864 40186 35873
rect 34426 35799 34482 35808
rect 35716 35828 35768 35834
rect 33140 35770 33192 35776
rect 35716 35770 35768 35776
rect 40040 35828 40092 35834
rect 40130 35799 40186 35808
rect 40040 35770 40092 35776
rect 31576 35760 31628 35766
rect 29092 35702 29144 35708
rect 30010 35728 30066 35737
rect 23570 35663 23626 35672
rect 30010 35663 30066 35672
rect 31022 35728 31078 35737
rect 33152 35737 33180 35770
rect 33600 35760 33652 35766
rect 31576 35702 31628 35708
rect 33138 35728 33194 35737
rect 31022 35663 31078 35672
rect 33138 35663 33194 35672
rect 33598 35728 33600 35737
rect 40052 35737 40080 35770
rect 42720 35737 42748 36343
rect 44088 36304 44140 36310
rect 44088 36246 44140 36252
rect 43536 36168 43588 36174
rect 43536 36110 43588 36116
rect 43548 35873 43576 36110
rect 44100 35902 44128 36246
rect 44088 35896 44140 35902
rect 43534 35864 43590 35873
rect 44088 35838 44140 35844
rect 43534 35799 43590 35808
rect 56060 35737 56088 37266
rect 56244 37262 56272 37810
rect 56612 37262 56640 40938
rect 56704 39370 56732 41006
rect 56784 39432 56836 39438
rect 56784 39374 56836 39380
rect 56692 39364 56744 39370
rect 56692 39306 56744 39312
rect 56796 38758 56824 39374
rect 57440 38962 57468 41006
rect 59280 39574 59308 42298
rect 59268 39568 59320 39574
rect 59268 39510 59320 39516
rect 59176 39296 59228 39302
rect 59176 39238 59228 39244
rect 59188 38962 59216 39238
rect 57428 38956 57480 38962
rect 57428 38898 57480 38904
rect 59176 38956 59228 38962
rect 59176 38898 59228 38904
rect 57796 38888 57848 38894
rect 57796 38830 57848 38836
rect 56784 38752 56836 38758
rect 56784 38694 56836 38700
rect 56690 37904 56746 37913
rect 56690 37839 56746 37848
rect 56704 37618 56732 37839
rect 56796 37738 56824 38694
rect 56876 38344 56928 38350
rect 56876 38286 56928 38292
rect 57152 38344 57204 38350
rect 57152 38286 57204 38292
rect 57704 38344 57756 38350
rect 57704 38286 57756 38292
rect 56888 37942 56916 38286
rect 57164 38010 57192 38286
rect 57716 38214 57744 38286
rect 57704 38208 57756 38214
rect 57704 38150 57756 38156
rect 57808 38010 57836 38830
rect 58164 38752 58216 38758
rect 58164 38694 58216 38700
rect 59176 38752 59228 38758
rect 59176 38694 59228 38700
rect 57152 38004 57204 38010
rect 57152 37946 57204 37952
rect 57796 38004 57848 38010
rect 57796 37946 57848 37952
rect 56876 37936 56928 37942
rect 56876 37878 56928 37884
rect 56784 37732 56836 37738
rect 56784 37674 56836 37680
rect 56876 37732 56928 37738
rect 56876 37674 56928 37680
rect 56888 37618 56916 37674
rect 56704 37590 56916 37618
rect 56704 37466 56732 37590
rect 56692 37460 56744 37466
rect 56692 37402 56744 37408
rect 57164 37330 57192 37946
rect 58176 37874 58204 38694
rect 59188 38214 59216 38694
rect 59280 38486 59308 39510
rect 59912 39364 59964 39370
rect 59912 39306 59964 39312
rect 59544 39024 59596 39030
rect 59544 38966 59596 38972
rect 59556 38486 59584 38966
rect 59636 38956 59688 38962
rect 59636 38898 59688 38904
rect 59268 38480 59320 38486
rect 59268 38422 59320 38428
rect 59544 38480 59596 38486
rect 59544 38422 59596 38428
rect 59176 38208 59228 38214
rect 59176 38150 59228 38156
rect 58164 37868 58216 37874
rect 58164 37810 58216 37816
rect 58256 37868 58308 37874
rect 58256 37810 58308 37816
rect 58268 37738 58296 37810
rect 59280 37806 59308 38422
rect 59268 37800 59320 37806
rect 59004 37748 59268 37754
rect 59004 37742 59320 37748
rect 58256 37732 58308 37738
rect 58256 37674 58308 37680
rect 59004 37726 59308 37742
rect 58072 37664 58124 37670
rect 58072 37606 58124 37612
rect 58084 37466 58112 37606
rect 58072 37460 58124 37466
rect 58072 37402 58124 37408
rect 59004 37330 59032 37726
rect 59280 37466 59308 37726
rect 59648 37670 59676 38898
rect 59924 38214 59952 39306
rect 60280 39296 60332 39302
rect 60280 39238 60332 39244
rect 60372 39296 60424 39302
rect 60372 39238 60424 39244
rect 60292 38894 60320 39238
rect 60280 38888 60332 38894
rect 60280 38830 60332 38836
rect 60384 38554 60412 39238
rect 60464 39092 60516 39098
rect 60464 39034 60516 39040
rect 60476 38654 60504 39034
rect 60476 38626 60596 38654
rect 60004 38548 60056 38554
rect 60004 38490 60056 38496
rect 60372 38548 60424 38554
rect 60372 38490 60424 38496
rect 60016 38214 60044 38490
rect 60568 38350 60596 38626
rect 60372 38344 60424 38350
rect 60372 38286 60424 38292
rect 60556 38344 60608 38350
rect 60556 38286 60608 38292
rect 60280 38276 60332 38282
rect 60280 38218 60332 38224
rect 59912 38208 59964 38214
rect 59912 38150 59964 38156
rect 60004 38208 60056 38214
rect 60004 38150 60056 38156
rect 60292 37806 60320 38218
rect 60384 38010 60412 38286
rect 60372 38004 60424 38010
rect 60372 37946 60424 37952
rect 60280 37800 60332 37806
rect 60280 37742 60332 37748
rect 59636 37664 59688 37670
rect 59636 37606 59688 37612
rect 59820 37664 59872 37670
rect 59820 37606 59872 37612
rect 59268 37460 59320 37466
rect 59268 37402 59320 37408
rect 59832 37398 59860 37606
rect 59820 37392 59872 37398
rect 59820 37334 59872 37340
rect 57152 37324 57204 37330
rect 57152 37266 57204 37272
rect 58992 37324 59044 37330
rect 58992 37266 59044 37272
rect 56232 37256 56284 37262
rect 56232 37198 56284 37204
rect 56600 37256 56652 37262
rect 56600 37198 56652 37204
rect 60568 35834 60596 38286
rect 60660 36786 60688 43046
rect 62672 42288 62724 42294
rect 62672 42230 62724 42236
rect 60738 41576 60794 41585
rect 60738 41511 60794 41520
rect 60752 40118 60780 41511
rect 62684 41414 62712 42230
rect 63040 42152 63092 42158
rect 63040 42094 63092 42100
rect 62684 41386 62988 41414
rect 60740 40112 60792 40118
rect 60740 40054 60792 40060
rect 62670 40080 62726 40089
rect 62670 40015 62726 40024
rect 62488 37800 62540 37806
rect 62488 37742 62540 37748
rect 62500 37466 62528 37742
rect 62488 37460 62540 37466
rect 62488 37402 62540 37408
rect 62500 37330 62528 37402
rect 62488 37324 62540 37330
rect 62488 37266 62540 37272
rect 60648 36780 60700 36786
rect 60648 36722 60700 36728
rect 61568 36304 61620 36310
rect 61568 36246 61620 36252
rect 60556 35828 60608 35834
rect 60556 35770 60608 35776
rect 33652 35728 33654 35737
rect 33598 35663 33654 35672
rect 40038 35728 40094 35737
rect 40038 35663 40094 35672
rect 42706 35728 42762 35737
rect 42706 35663 42762 35672
rect 56046 35728 56102 35737
rect 56046 35663 56102 35672
rect 22204 35562 22232 35663
rect 61580 35630 61608 36246
rect 62580 36032 62632 36038
rect 62580 35974 62632 35980
rect 61568 35624 61620 35630
rect 61568 35566 61620 35572
rect 62488 35624 62540 35630
rect 62488 35566 62540 35572
rect 8208 35556 8260 35562
rect 8208 35498 8260 35504
rect 18052 35556 18104 35562
rect 18052 35498 18104 35504
rect 22192 35556 22244 35562
rect 22192 35498 22244 35504
rect 62500 26234 62528 35566
rect 62592 35057 62620 35974
rect 62578 35048 62634 35057
rect 62578 34983 62634 34992
rect 62684 31754 62712 40015
rect 62856 36916 62908 36922
rect 62856 36858 62908 36864
rect 62762 36272 62818 36281
rect 62762 36207 62818 36216
rect 62592 31726 62712 31754
rect 62592 30924 62620 31726
rect 62670 30938 62726 30947
rect 62592 30896 62670 30924
rect 62670 30873 62726 30882
rect 62776 29247 62804 36207
rect 62762 29238 62818 29247
rect 62762 29173 62818 29182
rect 62500 26206 62804 26234
rect 62578 17232 62634 17241
rect 62578 17167 62634 17176
rect 62592 6914 62620 17167
rect 62500 6886 62620 6914
rect 48964 2032 49016 2038
rect 48964 1974 49016 1980
rect 48976 1873 49004 1974
rect 62500 1970 62528 6886
rect 49608 1964 49660 1970
rect 49608 1906 49660 1912
rect 62488 1964 62540 1970
rect 62488 1906 62540 1912
rect 49620 1873 49648 1906
rect 49700 1896 49752 1902
rect 48962 1864 49018 1873
rect 48962 1799 49018 1808
rect 49606 1864 49662 1873
rect 49700 1838 49752 1844
rect 49606 1799 49662 1808
rect 49712 1737 49740 1838
rect 49698 1728 49754 1737
rect 49698 1663 49754 1672
rect 62776 1465 62804 26206
rect 62868 6866 62896 36858
rect 62960 35290 62988 41386
rect 62948 35284 63000 35290
rect 62948 35226 63000 35232
rect 62960 34610 62988 35226
rect 62948 34604 63000 34610
rect 62948 34546 63000 34552
rect 62948 29980 63000 29986
rect 62948 29922 63000 29928
rect 62960 16726 62988 29922
rect 63052 23526 63080 42094
rect 63590 41168 63646 41177
rect 63590 41103 63646 41112
rect 64880 41132 64932 41138
rect 63500 39636 63552 39642
rect 63500 39578 63552 39584
rect 63132 38208 63184 38214
rect 63132 38150 63184 38156
rect 63144 29986 63172 38150
rect 63408 37800 63460 37806
rect 63408 37742 63460 37748
rect 63314 36544 63370 36553
rect 63314 36479 63370 36488
rect 63224 36304 63276 36310
rect 63224 36246 63276 36252
rect 63236 33998 63264 36246
rect 63224 33992 63276 33998
rect 63224 33934 63276 33940
rect 63132 29980 63184 29986
rect 63132 29922 63184 29928
rect 63328 28762 63356 36479
rect 63420 34134 63448 37742
rect 63512 36310 63540 39578
rect 63500 36304 63552 36310
rect 63500 36246 63552 36252
rect 63498 36136 63554 36145
rect 63498 36071 63554 36080
rect 63408 34128 63460 34134
rect 63408 34070 63460 34076
rect 63512 33153 63540 36071
rect 63604 35698 63632 41103
rect 64880 41074 64932 41080
rect 64694 39400 64750 39409
rect 64694 39335 64750 39344
rect 64236 38412 64288 38418
rect 64236 38354 64288 38360
rect 63960 37868 64012 37874
rect 63960 37810 64012 37816
rect 63868 37256 63920 37262
rect 63868 37198 63920 37204
rect 63880 36922 63908 37198
rect 63868 36916 63920 36922
rect 63868 36858 63920 36864
rect 63684 36236 63736 36242
rect 63684 36178 63736 36184
rect 63592 35692 63644 35698
rect 63592 35634 63644 35640
rect 63590 35592 63646 35601
rect 63590 35527 63646 35536
rect 63498 33144 63554 33153
rect 63498 33079 63554 33088
rect 63604 32994 63632 35527
rect 63696 34406 63724 36178
rect 63776 36168 63828 36174
rect 63776 36110 63828 36116
rect 63868 36168 63920 36174
rect 63868 36110 63920 36116
rect 63788 36009 63816 36110
rect 63774 36000 63830 36009
rect 63774 35935 63830 35944
rect 63880 35737 63908 36110
rect 63972 35766 64000 37810
rect 64052 37664 64104 37670
rect 64052 37606 64104 37612
rect 64064 36718 64092 37606
rect 64248 37330 64276 38354
rect 64236 37324 64288 37330
rect 64236 37266 64288 37272
rect 64052 36712 64104 36718
rect 64052 36654 64104 36660
rect 64144 36576 64196 36582
rect 64144 36518 64196 36524
rect 64156 36310 64184 36518
rect 64144 36304 64196 36310
rect 64144 36246 64196 36252
rect 63960 35760 64012 35766
rect 63866 35728 63922 35737
rect 63960 35702 64012 35708
rect 63866 35663 63922 35672
rect 63776 35624 63828 35630
rect 63776 35566 63828 35572
rect 63684 34400 63736 34406
rect 63684 34342 63736 34348
rect 63788 33946 63816 35566
rect 63880 35086 63908 35663
rect 63960 35624 64012 35630
rect 63960 35566 64012 35572
rect 63868 35080 63920 35086
rect 63868 35022 63920 35028
rect 63972 34202 64000 35566
rect 64052 35556 64104 35562
rect 64052 35498 64104 35504
rect 64064 34474 64092 35498
rect 64144 35488 64196 35494
rect 64144 35430 64196 35436
rect 64156 35222 64184 35430
rect 64144 35216 64196 35222
rect 64144 35158 64196 35164
rect 64144 35080 64196 35086
rect 64144 35022 64196 35028
rect 64052 34468 64104 34474
rect 64052 34410 64104 34416
rect 63960 34196 64012 34202
rect 63960 34138 64012 34144
rect 64156 34082 64184 35022
rect 63512 32966 63632 32994
rect 63696 33918 63816 33946
rect 63972 34054 64184 34082
rect 63512 31754 63540 32966
rect 63420 31726 63540 31754
rect 63316 28756 63368 28762
rect 63316 28698 63368 28704
rect 63328 28218 63356 28698
rect 63316 28212 63368 28218
rect 63316 28154 63368 28160
rect 63224 24880 63276 24886
rect 63224 24822 63276 24828
rect 63040 23520 63092 23526
rect 63040 23462 63092 23468
rect 63040 18420 63092 18426
rect 63040 18362 63092 18368
rect 62948 16720 63000 16726
rect 62948 16662 63000 16668
rect 62948 11688 63000 11694
rect 62948 11630 63000 11636
rect 62856 6860 62908 6866
rect 62856 6802 62908 6808
rect 62762 1456 62818 1465
rect 62762 1391 62818 1400
rect 62960 1329 62988 11630
rect 63052 2038 63080 18362
rect 63236 9654 63264 24822
rect 63316 21412 63368 21418
rect 63316 21354 63368 21360
rect 63328 16658 63356 21354
rect 63420 18034 63448 31726
rect 63696 28994 63724 33918
rect 63776 33856 63828 33862
rect 63776 33798 63828 33804
rect 63604 28966 63724 28994
rect 63604 24886 63632 28966
rect 63788 26234 63816 33798
rect 63868 30796 63920 30802
rect 63868 30738 63920 30744
rect 63880 26246 63908 30738
rect 63696 26206 63816 26234
rect 63868 26240 63920 26246
rect 63592 24880 63644 24886
rect 63592 24822 63644 24828
rect 63420 18006 63540 18034
rect 63316 16652 63368 16658
rect 63316 16594 63368 16600
rect 63512 16538 63540 18006
rect 63328 16510 63540 16538
rect 63224 9648 63276 9654
rect 63224 9590 63276 9596
rect 63328 6914 63356 16510
rect 63500 16448 63552 16454
rect 63500 16390 63552 16396
rect 63512 8974 63540 16390
rect 63500 8968 63552 8974
rect 63500 8910 63552 8916
rect 63328 6886 63540 6914
rect 63512 3670 63540 6886
rect 63592 6860 63644 6866
rect 63592 6802 63644 6808
rect 63604 5914 63632 6802
rect 63592 5908 63644 5914
rect 63592 5850 63644 5856
rect 63592 5772 63644 5778
rect 63592 5714 63644 5720
rect 63500 3664 63552 3670
rect 63500 3606 63552 3612
rect 63604 2650 63632 5714
rect 63592 2644 63644 2650
rect 63592 2586 63644 2592
rect 63040 2032 63092 2038
rect 63040 1974 63092 1980
rect 63696 1873 63724 26206
rect 63868 26182 63920 26188
rect 63972 25650 64000 34054
rect 64144 33992 64196 33998
rect 64144 33934 64196 33940
rect 64052 32972 64104 32978
rect 64052 32914 64104 32920
rect 64064 31482 64092 32914
rect 64156 31754 64184 33934
rect 64248 33046 64276 37266
rect 64338 37020 64646 37029
rect 64338 37018 64344 37020
rect 64400 37018 64424 37020
rect 64480 37018 64504 37020
rect 64560 37018 64584 37020
rect 64640 37018 64646 37020
rect 64400 36966 64402 37018
rect 64582 36966 64584 37018
rect 64338 36964 64344 36966
rect 64400 36964 64424 36966
rect 64480 36964 64504 36966
rect 64560 36964 64584 36966
rect 64640 36964 64646 36966
rect 64338 36955 64646 36964
rect 64338 35932 64646 35941
rect 64338 35930 64344 35932
rect 64400 35930 64424 35932
rect 64480 35930 64504 35932
rect 64560 35930 64584 35932
rect 64640 35930 64646 35932
rect 64400 35878 64402 35930
rect 64582 35878 64584 35930
rect 64338 35876 64344 35878
rect 64400 35876 64424 35878
rect 64480 35876 64504 35878
rect 64560 35876 64584 35878
rect 64640 35876 64646 35878
rect 64338 35867 64646 35876
rect 64708 35714 64736 39335
rect 64788 36644 64840 36650
rect 64788 36586 64840 36592
rect 64616 35686 64736 35714
rect 64616 35086 64644 35686
rect 64696 35488 64748 35494
rect 64696 35430 64748 35436
rect 64604 35080 64656 35086
rect 64604 35022 64656 35028
rect 64338 34844 64646 34853
rect 64338 34842 64344 34844
rect 64400 34842 64424 34844
rect 64480 34842 64504 34844
rect 64560 34842 64584 34844
rect 64640 34842 64646 34844
rect 64400 34790 64402 34842
rect 64582 34790 64584 34842
rect 64338 34788 64344 34790
rect 64400 34788 64424 34790
rect 64480 34788 64504 34790
rect 64560 34788 64584 34790
rect 64640 34788 64646 34790
rect 64338 34779 64646 34788
rect 64708 34746 64736 35430
rect 64696 34740 64748 34746
rect 64696 34682 64748 34688
rect 64800 34678 64828 36586
rect 64788 34672 64840 34678
rect 64788 34614 64840 34620
rect 64328 34468 64380 34474
rect 64328 34410 64380 34416
rect 64340 34134 64368 34410
rect 64788 34400 64840 34406
rect 64788 34342 64840 34348
rect 64328 34128 64380 34134
rect 64328 34070 64380 34076
rect 64338 33756 64646 33765
rect 64338 33754 64344 33756
rect 64400 33754 64424 33756
rect 64480 33754 64504 33756
rect 64560 33754 64584 33756
rect 64640 33754 64646 33756
rect 64400 33702 64402 33754
rect 64582 33702 64584 33754
rect 64338 33700 64344 33702
rect 64400 33700 64424 33702
rect 64480 33700 64504 33702
rect 64560 33700 64584 33702
rect 64640 33700 64646 33702
rect 64338 33691 64646 33700
rect 64328 33312 64380 33318
rect 64328 33254 64380 33260
rect 64340 33046 64368 33254
rect 64236 33040 64288 33046
rect 64236 32982 64288 32988
rect 64328 33040 64380 33046
rect 64328 32982 64380 32988
rect 64338 32668 64646 32677
rect 64338 32666 64344 32668
rect 64400 32666 64424 32668
rect 64480 32666 64504 32668
rect 64560 32666 64584 32668
rect 64640 32666 64646 32668
rect 64400 32614 64402 32666
rect 64582 32614 64584 32666
rect 64338 32612 64344 32614
rect 64400 32612 64424 32614
rect 64480 32612 64504 32614
rect 64560 32612 64584 32614
rect 64640 32612 64646 32614
rect 64338 32603 64646 32612
rect 64694 32464 64750 32473
rect 64694 32399 64750 32408
rect 64708 32366 64736 32399
rect 64696 32360 64748 32366
rect 64696 32302 64748 32308
rect 64156 31726 64276 31754
rect 64052 31476 64104 31482
rect 64052 31418 64104 31424
rect 64064 29170 64092 31418
rect 64052 29164 64104 29170
rect 64052 29106 64104 29112
rect 64052 26240 64104 26246
rect 64248 26234 64276 31726
rect 64338 31580 64646 31589
rect 64338 31578 64344 31580
rect 64400 31578 64424 31580
rect 64480 31578 64504 31580
rect 64560 31578 64584 31580
rect 64640 31578 64646 31580
rect 64400 31526 64402 31578
rect 64582 31526 64584 31578
rect 64338 31524 64344 31526
rect 64400 31524 64424 31526
rect 64480 31524 64504 31526
rect 64560 31524 64584 31526
rect 64640 31524 64646 31526
rect 64338 31515 64646 31524
rect 64338 30492 64646 30501
rect 64338 30490 64344 30492
rect 64400 30490 64424 30492
rect 64480 30490 64504 30492
rect 64560 30490 64584 30492
rect 64640 30490 64646 30492
rect 64400 30438 64402 30490
rect 64582 30438 64584 30490
rect 64338 30436 64344 30438
rect 64400 30436 64424 30438
rect 64480 30436 64504 30438
rect 64560 30436 64584 30438
rect 64640 30436 64646 30438
rect 64338 30427 64646 30436
rect 64328 30116 64380 30122
rect 64328 30058 64380 30064
rect 64340 29850 64368 30058
rect 64328 29844 64380 29850
rect 64328 29786 64380 29792
rect 64696 29504 64748 29510
rect 64696 29446 64748 29452
rect 64338 29404 64646 29413
rect 64338 29402 64344 29404
rect 64400 29402 64424 29404
rect 64480 29402 64504 29404
rect 64560 29402 64584 29404
rect 64640 29402 64646 29404
rect 64400 29350 64402 29402
rect 64582 29350 64584 29402
rect 64338 29348 64344 29350
rect 64400 29348 64424 29350
rect 64480 29348 64504 29350
rect 64560 29348 64584 29350
rect 64640 29348 64646 29350
rect 64338 29339 64646 29348
rect 64708 29170 64736 29446
rect 64696 29164 64748 29170
rect 64696 29106 64748 29112
rect 64338 28316 64646 28325
rect 64338 28314 64344 28316
rect 64400 28314 64424 28316
rect 64480 28314 64504 28316
rect 64560 28314 64584 28316
rect 64640 28314 64646 28316
rect 64400 28262 64402 28314
rect 64582 28262 64584 28314
rect 64338 28260 64344 28262
rect 64400 28260 64424 28262
rect 64480 28260 64504 28262
rect 64560 28260 64584 28262
rect 64640 28260 64646 28262
rect 64338 28251 64646 28260
rect 64338 27228 64646 27237
rect 64338 27226 64344 27228
rect 64400 27226 64424 27228
rect 64480 27226 64504 27228
rect 64560 27226 64584 27228
rect 64640 27226 64646 27228
rect 64400 27174 64402 27226
rect 64582 27174 64584 27226
rect 64338 27172 64344 27174
rect 64400 27172 64424 27174
rect 64480 27172 64504 27174
rect 64560 27172 64584 27174
rect 64640 27172 64646 27174
rect 64338 27163 64646 27172
rect 64696 26988 64748 26994
rect 64696 26930 64748 26936
rect 64604 26852 64656 26858
rect 64604 26794 64656 26800
rect 64616 26586 64644 26794
rect 64604 26580 64656 26586
rect 64604 26522 64656 26528
rect 64052 26182 64104 26188
rect 64156 26206 64276 26234
rect 63788 25622 64000 25650
rect 63788 1902 63816 25622
rect 63960 25356 64012 25362
rect 63960 25298 64012 25304
rect 63972 24614 64000 25298
rect 63960 24608 64012 24614
rect 63960 24550 64012 24556
rect 63972 23662 64000 24550
rect 64064 24342 64092 26182
rect 64052 24336 64104 24342
rect 64052 24278 64104 24284
rect 63960 23656 64012 23662
rect 63960 23598 64012 23604
rect 63868 23520 63920 23526
rect 63868 23462 63920 23468
rect 63880 21418 63908 23462
rect 63972 22098 64000 23598
rect 64052 22568 64104 22574
rect 64052 22510 64104 22516
rect 63960 22092 64012 22098
rect 63960 22034 64012 22040
rect 63868 21412 63920 21418
rect 63868 21354 63920 21360
rect 63972 16114 64000 22034
rect 64064 19854 64092 22510
rect 64156 22506 64184 26206
rect 64338 26140 64646 26149
rect 64338 26138 64344 26140
rect 64400 26138 64424 26140
rect 64480 26138 64504 26140
rect 64560 26138 64584 26140
rect 64640 26138 64646 26140
rect 64400 26086 64402 26138
rect 64582 26086 64584 26138
rect 64338 26084 64344 26086
rect 64400 26084 64424 26086
rect 64480 26084 64504 26086
rect 64560 26084 64584 26086
rect 64640 26084 64646 26086
rect 64338 26075 64646 26084
rect 64236 25152 64288 25158
rect 64236 25094 64288 25100
rect 64248 23594 64276 25094
rect 64338 25052 64646 25061
rect 64338 25050 64344 25052
rect 64400 25050 64424 25052
rect 64480 25050 64504 25052
rect 64560 25050 64584 25052
rect 64640 25050 64646 25052
rect 64400 24998 64402 25050
rect 64582 24998 64584 25050
rect 64338 24996 64344 24998
rect 64400 24996 64424 24998
rect 64480 24996 64504 24998
rect 64560 24996 64584 24998
rect 64640 24996 64646 24998
rect 64338 24987 64646 24996
rect 64708 24410 64736 26930
rect 64696 24404 64748 24410
rect 64696 24346 64748 24352
rect 64338 23964 64646 23973
rect 64338 23962 64344 23964
rect 64400 23962 64424 23964
rect 64480 23962 64504 23964
rect 64560 23962 64584 23964
rect 64640 23962 64646 23964
rect 64400 23910 64402 23962
rect 64582 23910 64584 23962
rect 64338 23908 64344 23910
rect 64400 23908 64424 23910
rect 64480 23908 64504 23910
rect 64560 23908 64584 23910
rect 64640 23908 64646 23910
rect 64338 23899 64646 23908
rect 64236 23588 64288 23594
rect 64236 23530 64288 23536
rect 64338 22876 64646 22885
rect 64338 22874 64344 22876
rect 64400 22874 64424 22876
rect 64480 22874 64504 22876
rect 64560 22874 64584 22876
rect 64640 22874 64646 22876
rect 64400 22822 64402 22874
rect 64582 22822 64584 22874
rect 64338 22820 64344 22822
rect 64400 22820 64424 22822
rect 64480 22820 64504 22822
rect 64560 22820 64584 22822
rect 64640 22820 64646 22822
rect 64338 22811 64646 22820
rect 64708 22574 64736 24346
rect 64696 22568 64748 22574
rect 64696 22510 64748 22516
rect 64144 22500 64196 22506
rect 64144 22442 64196 22448
rect 64800 22094 64828 34342
rect 64892 30802 64920 41074
rect 65064 40724 65116 40730
rect 65064 40666 65116 40672
rect 64972 40112 65024 40118
rect 64972 40054 65024 40060
rect 64984 33862 65012 40054
rect 64972 33856 65024 33862
rect 64972 33798 65024 33804
rect 64972 33312 65024 33318
rect 64972 33254 65024 33260
rect 64984 32570 65012 33254
rect 64972 32564 65024 32570
rect 64972 32506 65024 32512
rect 64972 32224 65024 32230
rect 64972 32166 65024 32172
rect 64984 31890 65012 32166
rect 64972 31884 65024 31890
rect 64972 31826 65024 31832
rect 64970 31784 65026 31793
rect 64970 31719 64972 31728
rect 65024 31719 65026 31728
rect 64972 31690 65024 31696
rect 65076 31362 65104 40666
rect 65258 37564 65566 37573
rect 65258 37562 65264 37564
rect 65320 37562 65344 37564
rect 65400 37562 65424 37564
rect 65480 37562 65504 37564
rect 65560 37562 65566 37564
rect 65320 37510 65322 37562
rect 65502 37510 65504 37562
rect 65258 37508 65264 37510
rect 65320 37508 65344 37510
rect 65400 37508 65424 37510
rect 65480 37508 65504 37510
rect 65560 37508 65566 37510
rect 65258 37499 65566 37508
rect 65800 37460 65852 37466
rect 65800 37402 65852 37408
rect 65708 37256 65760 37262
rect 65708 37198 65760 37204
rect 65432 37120 65484 37126
rect 65432 37062 65484 37068
rect 65444 36718 65472 37062
rect 65432 36712 65484 36718
rect 65432 36654 65484 36660
rect 65614 36680 65670 36689
rect 65614 36615 65670 36624
rect 65156 36576 65208 36582
rect 65156 36518 65208 36524
rect 65168 35834 65196 36518
rect 65258 36476 65566 36485
rect 65258 36474 65264 36476
rect 65320 36474 65344 36476
rect 65400 36474 65424 36476
rect 65480 36474 65504 36476
rect 65560 36474 65566 36476
rect 65320 36422 65322 36474
rect 65502 36422 65504 36474
rect 65258 36420 65264 36422
rect 65320 36420 65344 36422
rect 65400 36420 65424 36422
rect 65480 36420 65504 36422
rect 65560 36420 65566 36422
rect 65258 36411 65566 36420
rect 65628 36122 65656 36615
rect 65536 36094 65656 36122
rect 65156 35828 65208 35834
rect 65156 35770 65208 35776
rect 65536 35698 65564 36094
rect 65720 36038 65748 37198
rect 65812 36310 65840 37402
rect 66168 36848 66220 36854
rect 66168 36790 66220 36796
rect 66076 36372 66128 36378
rect 66076 36314 66128 36320
rect 65800 36304 65852 36310
rect 65800 36246 65852 36252
rect 65708 36032 65760 36038
rect 65708 35974 65760 35980
rect 65156 35692 65208 35698
rect 65156 35634 65208 35640
rect 65524 35692 65576 35698
rect 65524 35634 65576 35640
rect 65616 35692 65668 35698
rect 65616 35634 65668 35640
rect 65168 35272 65196 35634
rect 65258 35388 65566 35397
rect 65258 35386 65264 35388
rect 65320 35386 65344 35388
rect 65400 35386 65424 35388
rect 65480 35386 65504 35388
rect 65560 35386 65566 35388
rect 65320 35334 65322 35386
rect 65502 35334 65504 35386
rect 65258 35332 65264 35334
rect 65320 35332 65344 35334
rect 65400 35332 65424 35334
rect 65480 35332 65504 35334
rect 65560 35332 65566 35334
rect 65258 35323 65566 35332
rect 65628 35290 65656 35634
rect 65616 35284 65668 35290
rect 65168 35244 65288 35272
rect 65156 34944 65208 34950
rect 65156 34886 65208 34892
rect 64984 31334 65104 31362
rect 64984 31278 65012 31334
rect 64972 31272 65024 31278
rect 64972 31214 65024 31220
rect 65064 31272 65116 31278
rect 65064 31214 65116 31220
rect 64880 30796 64932 30802
rect 64880 30738 64932 30744
rect 64880 30660 64932 30666
rect 64880 30602 64932 30608
rect 64892 28490 64920 30602
rect 64880 28484 64932 28490
rect 64880 28426 64932 28432
rect 64880 27532 64932 27538
rect 64880 27474 64932 27480
rect 64892 26314 64920 27474
rect 64880 26308 64932 26314
rect 64880 26250 64932 26256
rect 64984 24750 65012 31214
rect 65076 30666 65104 31214
rect 65168 30938 65196 34886
rect 65260 34610 65288 35244
rect 65616 35226 65668 35232
rect 65616 34944 65668 34950
rect 65616 34886 65668 34892
rect 65248 34604 65300 34610
rect 65248 34546 65300 34552
rect 65628 34542 65656 34886
rect 65616 34536 65668 34542
rect 65616 34478 65668 34484
rect 65258 34300 65566 34309
rect 65258 34298 65264 34300
rect 65320 34298 65344 34300
rect 65400 34298 65424 34300
rect 65480 34298 65504 34300
rect 65560 34298 65566 34300
rect 65320 34246 65322 34298
rect 65502 34246 65504 34298
rect 65258 34244 65264 34246
rect 65320 34244 65344 34246
rect 65400 34244 65424 34246
rect 65480 34244 65504 34246
rect 65560 34244 65566 34246
rect 65258 34235 65566 34244
rect 65628 34066 65656 34478
rect 65616 34060 65668 34066
rect 65616 34002 65668 34008
rect 65258 33212 65566 33221
rect 65258 33210 65264 33212
rect 65320 33210 65344 33212
rect 65400 33210 65424 33212
rect 65480 33210 65504 33212
rect 65560 33210 65566 33212
rect 65320 33158 65322 33210
rect 65502 33158 65504 33210
rect 65258 33156 65264 33158
rect 65320 33156 65344 33158
rect 65400 33156 65424 33158
rect 65480 33156 65504 33158
rect 65560 33156 65566 33158
rect 65258 33147 65566 33156
rect 65720 32434 65748 35974
rect 65812 35222 65840 36246
rect 65984 35556 66036 35562
rect 65984 35498 66036 35504
rect 65892 35284 65944 35290
rect 65892 35226 65944 35232
rect 65800 35216 65852 35222
rect 65800 35158 65852 35164
rect 65904 32502 65932 35226
rect 65996 33522 66024 35498
rect 65984 33516 66036 33522
rect 65984 33458 66036 33464
rect 65996 33114 66024 33458
rect 65984 33108 66036 33114
rect 65984 33050 66036 33056
rect 65892 32496 65944 32502
rect 65892 32438 65944 32444
rect 65708 32428 65760 32434
rect 65708 32370 65760 32376
rect 65258 32124 65566 32133
rect 65258 32122 65264 32124
rect 65320 32122 65344 32124
rect 65400 32122 65424 32124
rect 65480 32122 65504 32124
rect 65560 32122 65566 32124
rect 65320 32070 65322 32122
rect 65502 32070 65504 32122
rect 65258 32068 65264 32070
rect 65320 32068 65344 32070
rect 65400 32068 65424 32070
rect 65480 32068 65504 32070
rect 65560 32068 65566 32070
rect 65258 32059 65566 32068
rect 65800 32020 65852 32026
rect 65800 31962 65852 31968
rect 65616 31952 65668 31958
rect 65616 31894 65668 31900
rect 65340 31884 65392 31890
rect 65340 31826 65392 31832
rect 65248 31816 65300 31822
rect 65352 31793 65380 31826
rect 65248 31758 65300 31764
rect 65338 31784 65394 31793
rect 65260 31278 65288 31758
rect 65338 31719 65394 31728
rect 65248 31272 65300 31278
rect 65248 31214 65300 31220
rect 65258 31036 65566 31045
rect 65258 31034 65264 31036
rect 65320 31034 65344 31036
rect 65400 31034 65424 31036
rect 65480 31034 65504 31036
rect 65560 31034 65566 31036
rect 65320 30982 65322 31034
rect 65502 30982 65504 31034
rect 65258 30980 65264 30982
rect 65320 30980 65344 30982
rect 65400 30980 65424 30982
rect 65480 30980 65504 30982
rect 65560 30980 65566 30982
rect 65258 30971 65566 30980
rect 65156 30932 65208 30938
rect 65156 30874 65208 30880
rect 65064 30660 65116 30666
rect 65064 30602 65116 30608
rect 65168 30274 65196 30874
rect 65076 30258 65196 30274
rect 65064 30252 65196 30258
rect 65116 30246 65196 30252
rect 65064 30194 65116 30200
rect 65258 29948 65566 29957
rect 65258 29946 65264 29948
rect 65320 29946 65344 29948
rect 65400 29946 65424 29948
rect 65480 29946 65504 29948
rect 65560 29946 65566 29948
rect 65320 29894 65322 29946
rect 65502 29894 65504 29946
rect 65258 29892 65264 29894
rect 65320 29892 65344 29894
rect 65400 29892 65424 29894
rect 65480 29892 65504 29894
rect 65560 29892 65566 29894
rect 65258 29883 65566 29892
rect 65064 29776 65116 29782
rect 65064 29718 65116 29724
rect 65076 28694 65104 29718
rect 65156 29708 65208 29714
rect 65156 29650 65208 29656
rect 65168 28762 65196 29650
rect 65628 29306 65656 31894
rect 65708 31816 65760 31822
rect 65708 31758 65760 31764
rect 65720 29850 65748 31758
rect 65812 29850 65840 31962
rect 65904 31890 65932 32438
rect 65996 32230 66024 33050
rect 65984 32224 66036 32230
rect 65984 32166 66036 32172
rect 65892 31884 65944 31890
rect 65892 31826 65944 31832
rect 65890 31784 65946 31793
rect 65890 31719 65946 31728
rect 65984 31748 66036 31754
rect 65708 29844 65760 29850
rect 65708 29786 65760 29792
rect 65800 29844 65852 29850
rect 65800 29786 65852 29792
rect 65616 29300 65668 29306
rect 65616 29242 65668 29248
rect 65258 28860 65566 28869
rect 65258 28858 65264 28860
rect 65320 28858 65344 28860
rect 65400 28858 65424 28860
rect 65480 28858 65504 28860
rect 65560 28858 65566 28860
rect 65320 28806 65322 28858
rect 65502 28806 65504 28858
rect 65258 28804 65264 28806
rect 65320 28804 65344 28806
rect 65400 28804 65424 28806
rect 65480 28804 65504 28806
rect 65560 28804 65566 28806
rect 65258 28795 65566 28804
rect 65156 28756 65208 28762
rect 65156 28698 65208 28704
rect 65064 28688 65116 28694
rect 65064 28630 65116 28636
rect 65628 28626 65656 29242
rect 65800 29028 65852 29034
rect 65800 28970 65852 28976
rect 65616 28620 65668 28626
rect 65616 28562 65668 28568
rect 65156 28484 65208 28490
rect 65156 28426 65208 28432
rect 65168 27470 65196 28426
rect 65258 27772 65566 27781
rect 65258 27770 65264 27772
rect 65320 27770 65344 27772
rect 65400 27770 65424 27772
rect 65480 27770 65504 27772
rect 65560 27770 65566 27772
rect 65320 27718 65322 27770
rect 65502 27718 65504 27770
rect 65258 27716 65264 27718
rect 65320 27716 65344 27718
rect 65400 27716 65424 27718
rect 65480 27716 65504 27718
rect 65560 27716 65566 27718
rect 65258 27707 65566 27716
rect 65628 27674 65656 28562
rect 65616 27668 65668 27674
rect 65616 27610 65668 27616
rect 65156 27464 65208 27470
rect 65156 27406 65208 27412
rect 65708 27464 65760 27470
rect 65708 27406 65760 27412
rect 65064 27328 65116 27334
rect 65064 27270 65116 27276
rect 65076 26586 65104 27270
rect 65258 26684 65566 26693
rect 65258 26682 65264 26684
rect 65320 26682 65344 26684
rect 65400 26682 65424 26684
rect 65480 26682 65504 26684
rect 65560 26682 65566 26684
rect 65320 26630 65322 26682
rect 65502 26630 65504 26682
rect 65258 26628 65264 26630
rect 65320 26628 65344 26630
rect 65400 26628 65424 26630
rect 65480 26628 65504 26630
rect 65560 26628 65566 26630
rect 65258 26619 65566 26628
rect 65064 26580 65116 26586
rect 65064 26522 65116 26528
rect 65524 26580 65576 26586
rect 65524 26522 65576 26528
rect 65156 26376 65208 26382
rect 65156 26318 65208 26324
rect 65168 25294 65196 26318
rect 65536 26234 65564 26522
rect 65536 26206 65656 26234
rect 65258 25596 65566 25605
rect 65258 25594 65264 25596
rect 65320 25594 65344 25596
rect 65400 25594 65424 25596
rect 65480 25594 65504 25596
rect 65560 25594 65566 25596
rect 65320 25542 65322 25594
rect 65502 25542 65504 25594
rect 65258 25540 65264 25542
rect 65320 25540 65344 25542
rect 65400 25540 65424 25542
rect 65480 25540 65504 25542
rect 65560 25540 65566 25542
rect 65258 25531 65566 25540
rect 65064 25288 65116 25294
rect 65064 25230 65116 25236
rect 65156 25288 65208 25294
rect 65156 25230 65208 25236
rect 64972 24744 65024 24750
rect 64972 24686 65024 24692
rect 65076 23322 65104 25230
rect 65258 24508 65566 24517
rect 65258 24506 65264 24508
rect 65320 24506 65344 24508
rect 65400 24506 65424 24508
rect 65480 24506 65504 24508
rect 65560 24506 65566 24508
rect 65320 24454 65322 24506
rect 65502 24454 65504 24506
rect 65258 24452 65264 24454
rect 65320 24452 65344 24454
rect 65400 24452 65424 24454
rect 65480 24452 65504 24454
rect 65560 24452 65566 24454
rect 65258 24443 65566 24452
rect 65628 23594 65656 26206
rect 65616 23588 65668 23594
rect 65616 23530 65668 23536
rect 65258 23420 65566 23429
rect 65258 23418 65264 23420
rect 65320 23418 65344 23420
rect 65400 23418 65424 23420
rect 65480 23418 65504 23420
rect 65560 23418 65566 23420
rect 65320 23366 65322 23418
rect 65502 23366 65504 23418
rect 65258 23364 65264 23366
rect 65320 23364 65344 23366
rect 65400 23364 65424 23366
rect 65480 23364 65504 23366
rect 65560 23364 65566 23366
rect 65258 23355 65566 23364
rect 65064 23316 65116 23322
rect 65064 23258 65116 23264
rect 64880 23180 64932 23186
rect 64880 23122 64932 23128
rect 64892 22778 64920 23122
rect 65720 23118 65748 27406
rect 65812 26926 65840 28970
rect 65800 26920 65852 26926
rect 65800 26862 65852 26868
rect 65800 26784 65852 26790
rect 65800 26726 65852 26732
rect 65812 26450 65840 26726
rect 65800 26444 65852 26450
rect 65800 26386 65852 26392
rect 65800 26308 65852 26314
rect 65800 26250 65852 26256
rect 65812 25294 65840 26250
rect 65800 25288 65852 25294
rect 65800 25230 65852 25236
rect 65812 23526 65840 25230
rect 65800 23520 65852 23526
rect 65800 23462 65852 23468
rect 65708 23112 65760 23118
rect 65708 23054 65760 23060
rect 64880 22772 64932 22778
rect 64880 22714 64932 22720
rect 64880 22500 64932 22506
rect 64880 22442 64932 22448
rect 64248 22066 64828 22094
rect 64144 20324 64196 20330
rect 64144 20266 64196 20272
rect 64052 19848 64104 19854
rect 64052 19790 64104 19796
rect 64064 18222 64092 19790
rect 64052 18216 64104 18222
rect 64052 18158 64104 18164
rect 63960 16108 64012 16114
rect 63960 16050 64012 16056
rect 63972 12850 64000 16050
rect 63960 12844 64012 12850
rect 63960 12786 64012 12792
rect 63972 12434 64000 12786
rect 63880 12406 64000 12434
rect 63880 12238 63908 12406
rect 63868 12232 63920 12238
rect 63868 12174 63920 12180
rect 63880 10062 63908 12174
rect 63868 10056 63920 10062
rect 63868 9998 63920 10004
rect 63880 4690 63908 9998
rect 63960 9648 64012 9654
rect 63960 9590 64012 9596
rect 63972 6254 64000 9590
rect 64064 7954 64092 18158
rect 64156 11694 64184 20266
rect 64144 11688 64196 11694
rect 64144 11630 64196 11636
rect 64248 9058 64276 22066
rect 64696 22024 64748 22030
rect 64696 21966 64748 21972
rect 64338 21788 64646 21797
rect 64338 21786 64344 21788
rect 64400 21786 64424 21788
rect 64480 21786 64504 21788
rect 64560 21786 64584 21788
rect 64640 21786 64646 21788
rect 64400 21734 64402 21786
rect 64582 21734 64584 21786
rect 64338 21732 64344 21734
rect 64400 21732 64424 21734
rect 64480 21732 64504 21734
rect 64560 21732 64584 21734
rect 64640 21732 64646 21734
rect 64338 21723 64646 21732
rect 64708 21146 64736 21966
rect 64696 21140 64748 21146
rect 64696 21082 64748 21088
rect 64338 20700 64646 20709
rect 64338 20698 64344 20700
rect 64400 20698 64424 20700
rect 64480 20698 64504 20700
rect 64560 20698 64584 20700
rect 64640 20698 64646 20700
rect 64400 20646 64402 20698
rect 64582 20646 64584 20698
rect 64338 20644 64344 20646
rect 64400 20644 64424 20646
rect 64480 20644 64504 20646
rect 64560 20644 64584 20646
rect 64640 20644 64646 20646
rect 64338 20635 64646 20644
rect 64892 20346 64920 22442
rect 65258 22332 65566 22341
rect 65258 22330 65264 22332
rect 65320 22330 65344 22332
rect 65400 22330 65424 22332
rect 65480 22330 65504 22332
rect 65560 22330 65566 22332
rect 65320 22278 65322 22330
rect 65502 22278 65504 22330
rect 65258 22276 65264 22278
rect 65320 22276 65344 22278
rect 65400 22276 65424 22278
rect 65480 22276 65504 22278
rect 65560 22276 65566 22278
rect 65258 22267 65566 22276
rect 65708 21480 65760 21486
rect 65708 21422 65760 21428
rect 65616 21412 65668 21418
rect 65616 21354 65668 21360
rect 65156 21344 65208 21350
rect 65156 21286 65208 21292
rect 65168 21146 65196 21286
rect 65258 21244 65566 21253
rect 65258 21242 65264 21244
rect 65320 21242 65344 21244
rect 65400 21242 65424 21244
rect 65480 21242 65504 21244
rect 65560 21242 65566 21244
rect 65320 21190 65322 21242
rect 65502 21190 65504 21242
rect 65258 21188 65264 21190
rect 65320 21188 65344 21190
rect 65400 21188 65424 21190
rect 65480 21188 65504 21190
rect 65560 21188 65566 21190
rect 65258 21179 65566 21188
rect 65156 21140 65208 21146
rect 65156 21082 65208 21088
rect 65628 20942 65656 21354
rect 65064 20936 65116 20942
rect 65064 20878 65116 20884
rect 65616 20936 65668 20942
rect 65616 20878 65668 20884
rect 64972 20460 65024 20466
rect 64972 20402 65024 20408
rect 64800 20318 64920 20346
rect 64696 19848 64748 19854
rect 64696 19790 64748 19796
rect 64338 19612 64646 19621
rect 64338 19610 64344 19612
rect 64400 19610 64424 19612
rect 64480 19610 64504 19612
rect 64560 19610 64584 19612
rect 64640 19610 64646 19612
rect 64400 19558 64402 19610
rect 64582 19558 64584 19610
rect 64338 19556 64344 19558
rect 64400 19556 64424 19558
rect 64480 19556 64504 19558
rect 64560 19556 64584 19558
rect 64640 19556 64646 19558
rect 64338 19547 64646 19556
rect 64708 19514 64736 19790
rect 64696 19508 64748 19514
rect 64696 19450 64748 19456
rect 64696 18624 64748 18630
rect 64696 18566 64748 18572
rect 64338 18524 64646 18533
rect 64338 18522 64344 18524
rect 64400 18522 64424 18524
rect 64480 18522 64504 18524
rect 64560 18522 64584 18524
rect 64640 18522 64646 18524
rect 64400 18470 64402 18522
rect 64582 18470 64584 18522
rect 64338 18468 64344 18470
rect 64400 18468 64424 18470
rect 64480 18468 64504 18470
rect 64560 18468 64584 18470
rect 64640 18468 64646 18470
rect 64338 18459 64646 18468
rect 64708 18290 64736 18566
rect 64696 18284 64748 18290
rect 64696 18226 64748 18232
rect 64694 17912 64750 17921
rect 64694 17847 64750 17856
rect 64708 17814 64736 17847
rect 64696 17808 64748 17814
rect 64696 17750 64748 17756
rect 64338 17436 64646 17445
rect 64338 17434 64344 17436
rect 64400 17434 64424 17436
rect 64480 17434 64504 17436
rect 64560 17434 64584 17436
rect 64640 17434 64646 17436
rect 64400 17382 64402 17434
rect 64582 17382 64584 17434
rect 64338 17380 64344 17382
rect 64400 17380 64424 17382
rect 64480 17380 64504 17382
rect 64560 17380 64584 17382
rect 64640 17380 64646 17382
rect 64338 17371 64646 17380
rect 64708 17338 64736 17750
rect 64696 17332 64748 17338
rect 64696 17274 64748 17280
rect 64696 16448 64748 16454
rect 64696 16390 64748 16396
rect 64338 16348 64646 16357
rect 64338 16346 64344 16348
rect 64400 16346 64424 16348
rect 64480 16346 64504 16348
rect 64560 16346 64584 16348
rect 64640 16346 64646 16348
rect 64400 16294 64402 16346
rect 64582 16294 64584 16346
rect 64338 16292 64344 16294
rect 64400 16292 64424 16294
rect 64480 16292 64504 16294
rect 64560 16292 64584 16294
rect 64640 16292 64646 16294
rect 64338 16283 64646 16292
rect 64708 16114 64736 16390
rect 64696 16108 64748 16114
rect 64696 16050 64748 16056
rect 64800 15858 64828 20318
rect 64880 20256 64932 20262
rect 64880 20198 64932 20204
rect 64892 19310 64920 20198
rect 64880 19304 64932 19310
rect 64880 19246 64932 19252
rect 64984 19122 65012 20402
rect 64892 19094 65012 19122
rect 64892 17678 64920 19094
rect 65076 18850 65104 20878
rect 65258 20156 65566 20165
rect 65258 20154 65264 20156
rect 65320 20154 65344 20156
rect 65400 20154 65424 20156
rect 65480 20154 65504 20156
rect 65560 20154 65566 20156
rect 65320 20102 65322 20154
rect 65502 20102 65504 20154
rect 65258 20100 65264 20102
rect 65320 20100 65344 20102
rect 65400 20100 65424 20102
rect 65480 20100 65504 20102
rect 65560 20100 65566 20102
rect 65258 20091 65566 20100
rect 65628 19378 65656 20878
rect 65616 19372 65668 19378
rect 65616 19314 65668 19320
rect 65258 19068 65566 19077
rect 65258 19066 65264 19068
rect 65320 19066 65344 19068
rect 65400 19066 65424 19068
rect 65480 19066 65504 19068
rect 65560 19066 65566 19068
rect 65320 19014 65322 19066
rect 65502 19014 65504 19066
rect 65258 19012 65264 19014
rect 65320 19012 65344 19014
rect 65400 19012 65424 19014
rect 65480 19012 65504 19014
rect 65560 19012 65566 19014
rect 65258 19003 65566 19012
rect 65076 18822 65196 18850
rect 65064 18760 65116 18766
rect 65064 18702 65116 18708
rect 64972 18080 65024 18086
rect 64972 18022 65024 18028
rect 64984 17882 65012 18022
rect 65076 17882 65104 18702
rect 64972 17876 65024 17882
rect 64972 17818 65024 17824
rect 65064 17876 65116 17882
rect 65064 17818 65116 17824
rect 64880 17672 64932 17678
rect 64880 17614 64932 17620
rect 64708 15830 64828 15858
rect 64338 15260 64646 15269
rect 64338 15258 64344 15260
rect 64400 15258 64424 15260
rect 64480 15258 64504 15260
rect 64560 15258 64584 15260
rect 64640 15258 64646 15260
rect 64400 15206 64402 15258
rect 64582 15206 64584 15258
rect 64338 15204 64344 15206
rect 64400 15204 64424 15206
rect 64480 15204 64504 15206
rect 64560 15204 64584 15206
rect 64640 15204 64646 15206
rect 64338 15195 64646 15204
rect 64338 14172 64646 14181
rect 64338 14170 64344 14172
rect 64400 14170 64424 14172
rect 64480 14170 64504 14172
rect 64560 14170 64584 14172
rect 64640 14170 64646 14172
rect 64400 14118 64402 14170
rect 64582 14118 64584 14170
rect 64338 14116 64344 14118
rect 64400 14116 64424 14118
rect 64480 14116 64504 14118
rect 64560 14116 64584 14118
rect 64640 14116 64646 14118
rect 64338 14107 64646 14116
rect 64338 13084 64646 13093
rect 64338 13082 64344 13084
rect 64400 13082 64424 13084
rect 64480 13082 64504 13084
rect 64560 13082 64584 13084
rect 64640 13082 64646 13084
rect 64400 13030 64402 13082
rect 64582 13030 64584 13082
rect 64338 13028 64344 13030
rect 64400 13028 64424 13030
rect 64480 13028 64504 13030
rect 64560 13028 64584 13030
rect 64640 13028 64646 13030
rect 64338 13019 64646 13028
rect 64708 12730 64736 15830
rect 64786 15736 64842 15745
rect 64786 15671 64788 15680
rect 64840 15671 64842 15680
rect 64788 15642 64840 15648
rect 64800 15162 64828 15642
rect 64892 15502 64920 17614
rect 65168 17610 65196 18822
rect 65628 18766 65656 19314
rect 65616 18760 65668 18766
rect 65616 18702 65668 18708
rect 65258 17980 65566 17989
rect 65258 17978 65264 17980
rect 65320 17978 65344 17980
rect 65400 17978 65424 17980
rect 65480 17978 65504 17980
rect 65560 17978 65566 17980
rect 65320 17926 65322 17978
rect 65502 17926 65504 17978
rect 65258 17924 65264 17926
rect 65320 17924 65344 17926
rect 65400 17924 65424 17926
rect 65480 17924 65504 17926
rect 65560 17924 65566 17926
rect 65258 17915 65566 17924
rect 65156 17604 65208 17610
rect 65156 17546 65208 17552
rect 65258 16892 65566 16901
rect 65258 16890 65264 16892
rect 65320 16890 65344 16892
rect 65400 16890 65424 16892
rect 65480 16890 65504 16892
rect 65560 16890 65566 16892
rect 65320 16838 65322 16890
rect 65502 16838 65504 16890
rect 65258 16836 65264 16838
rect 65320 16836 65344 16838
rect 65400 16836 65424 16838
rect 65480 16836 65504 16838
rect 65560 16836 65566 16838
rect 65258 16827 65566 16836
rect 65064 16584 65116 16590
rect 65064 16526 65116 16532
rect 65076 15706 65104 16526
rect 65258 15804 65566 15813
rect 65258 15802 65264 15804
rect 65320 15802 65344 15804
rect 65400 15802 65424 15804
rect 65480 15802 65504 15804
rect 65560 15802 65566 15804
rect 65320 15750 65322 15802
rect 65502 15750 65504 15802
rect 65258 15748 65264 15750
rect 65320 15748 65344 15750
rect 65400 15748 65424 15750
rect 65480 15748 65504 15750
rect 65560 15748 65566 15750
rect 65258 15739 65566 15748
rect 65064 15700 65116 15706
rect 65064 15642 65116 15648
rect 64880 15496 64932 15502
rect 64880 15438 64932 15444
rect 65156 15496 65208 15502
rect 65156 15438 65208 15444
rect 64788 15156 64840 15162
rect 64788 15098 64840 15104
rect 65064 12844 65116 12850
rect 65064 12786 65116 12792
rect 64708 12714 64828 12730
rect 64708 12708 64840 12714
rect 64708 12702 64788 12708
rect 64788 12650 64840 12656
rect 64696 12232 64748 12238
rect 64696 12174 64748 12180
rect 64338 11996 64646 12005
rect 64338 11994 64344 11996
rect 64400 11994 64424 11996
rect 64480 11994 64504 11996
rect 64560 11994 64584 11996
rect 64640 11994 64646 11996
rect 64400 11942 64402 11994
rect 64582 11942 64584 11994
rect 64338 11940 64344 11942
rect 64400 11940 64424 11942
rect 64480 11940 64504 11942
rect 64560 11940 64584 11942
rect 64640 11940 64646 11942
rect 64338 11931 64646 11940
rect 64708 11898 64736 12174
rect 65076 11898 65104 12786
rect 64696 11892 64748 11898
rect 64696 11834 64748 11840
rect 65064 11892 65116 11898
rect 65064 11834 65116 11840
rect 64880 11552 64932 11558
rect 64880 11494 64932 11500
rect 64892 11354 64920 11494
rect 64880 11348 64932 11354
rect 64880 11290 64932 11296
rect 64338 10908 64646 10917
rect 64338 10906 64344 10908
rect 64400 10906 64424 10908
rect 64480 10906 64504 10908
rect 64560 10906 64584 10908
rect 64640 10906 64646 10908
rect 64400 10854 64402 10906
rect 64582 10854 64584 10906
rect 64338 10852 64344 10854
rect 64400 10852 64424 10854
rect 64480 10852 64504 10854
rect 64560 10852 64584 10854
rect 64640 10852 64646 10854
rect 64338 10843 64646 10852
rect 65168 10674 65196 15438
rect 65258 14716 65566 14725
rect 65258 14714 65264 14716
rect 65320 14714 65344 14716
rect 65400 14714 65424 14716
rect 65480 14714 65504 14716
rect 65560 14714 65566 14716
rect 65320 14662 65322 14714
rect 65502 14662 65504 14714
rect 65258 14660 65264 14662
rect 65320 14660 65344 14662
rect 65400 14660 65424 14662
rect 65480 14660 65504 14662
rect 65560 14660 65566 14662
rect 65258 14651 65566 14660
rect 65258 13628 65566 13637
rect 65258 13626 65264 13628
rect 65320 13626 65344 13628
rect 65400 13626 65424 13628
rect 65480 13626 65504 13628
rect 65560 13626 65566 13628
rect 65320 13574 65322 13626
rect 65502 13574 65504 13626
rect 65258 13572 65264 13574
rect 65320 13572 65344 13574
rect 65400 13572 65424 13574
rect 65480 13572 65504 13574
rect 65560 13572 65566 13574
rect 65258 13563 65566 13572
rect 65258 12540 65566 12549
rect 65258 12538 65264 12540
rect 65320 12538 65344 12540
rect 65400 12538 65424 12540
rect 65480 12538 65504 12540
rect 65560 12538 65566 12540
rect 65320 12486 65322 12538
rect 65502 12486 65504 12538
rect 65258 12484 65264 12486
rect 65320 12484 65344 12486
rect 65400 12484 65424 12486
rect 65480 12484 65504 12486
rect 65560 12484 65566 12486
rect 65258 12475 65566 12484
rect 65628 11762 65656 18702
rect 65720 17882 65748 21422
rect 65812 20398 65840 23462
rect 65904 23186 65932 31719
rect 65984 31690 66036 31696
rect 65996 30054 66024 31690
rect 65984 30048 66036 30054
rect 65984 29990 66036 29996
rect 65996 28762 66024 29990
rect 65984 28756 66036 28762
rect 65984 28698 66036 28704
rect 65984 26920 66036 26926
rect 65984 26862 66036 26868
rect 65996 26586 66024 26862
rect 65984 26580 66036 26586
rect 65984 26522 66036 26528
rect 65984 26444 66036 26450
rect 65984 26386 66036 26392
rect 65996 23254 66024 26386
rect 65984 23248 66036 23254
rect 65984 23190 66036 23196
rect 65892 23180 65944 23186
rect 65892 23122 65944 23128
rect 65892 22500 65944 22506
rect 65892 22442 65944 22448
rect 65904 22166 65932 22442
rect 65892 22160 65944 22166
rect 65892 22102 65944 22108
rect 65800 20392 65852 20398
rect 65800 20334 65852 20340
rect 65800 20256 65852 20262
rect 65800 20198 65852 20204
rect 65708 17876 65760 17882
rect 65708 17818 65760 17824
rect 65812 16658 65840 20198
rect 65904 19990 65932 22102
rect 65892 19984 65944 19990
rect 65892 19926 65944 19932
rect 65892 19712 65944 19718
rect 65892 19654 65944 19660
rect 65904 19310 65932 19654
rect 65892 19304 65944 19310
rect 65892 19246 65944 19252
rect 65800 16652 65852 16658
rect 65800 16594 65852 16600
rect 65812 16250 65840 16594
rect 65800 16244 65852 16250
rect 65800 16186 65852 16192
rect 65616 11756 65668 11762
rect 65616 11698 65668 11704
rect 65258 11452 65566 11461
rect 65258 11450 65264 11452
rect 65320 11450 65344 11452
rect 65400 11450 65424 11452
rect 65480 11450 65504 11452
rect 65560 11450 65566 11452
rect 65320 11398 65322 11450
rect 65502 11398 65504 11450
rect 65258 11396 65264 11398
rect 65320 11396 65344 11398
rect 65400 11396 65424 11398
rect 65480 11396 65504 11398
rect 65560 11396 65566 11398
rect 65258 11387 65566 11396
rect 65628 10826 65656 11698
rect 65628 10798 65748 10826
rect 65616 10736 65668 10742
rect 65616 10678 65668 10684
rect 65156 10668 65208 10674
rect 65156 10610 65208 10616
rect 64972 10464 65024 10470
rect 64972 10406 65024 10412
rect 64696 10056 64748 10062
rect 64696 9998 64748 10004
rect 64338 9820 64646 9829
rect 64338 9818 64344 9820
rect 64400 9818 64424 9820
rect 64480 9818 64504 9820
rect 64560 9818 64584 9820
rect 64640 9818 64646 9820
rect 64400 9766 64402 9818
rect 64582 9766 64584 9818
rect 64338 9764 64344 9766
rect 64400 9764 64424 9766
rect 64480 9764 64504 9766
rect 64560 9764 64584 9766
rect 64640 9764 64646 9766
rect 64338 9755 64646 9764
rect 64708 9178 64736 9998
rect 64984 9926 65012 10406
rect 64972 9920 65024 9926
rect 64972 9862 65024 9868
rect 64984 9518 65012 9862
rect 65168 9586 65196 10610
rect 65258 10364 65566 10373
rect 65258 10362 65264 10364
rect 65320 10362 65344 10364
rect 65400 10362 65424 10364
rect 65480 10362 65504 10364
rect 65560 10362 65566 10364
rect 65320 10310 65322 10362
rect 65502 10310 65504 10362
rect 65258 10308 65264 10310
rect 65320 10308 65344 10310
rect 65400 10308 65424 10310
rect 65480 10308 65504 10310
rect 65560 10308 65566 10310
rect 65258 10299 65566 10308
rect 65156 9580 65208 9586
rect 65156 9522 65208 9528
rect 64880 9512 64932 9518
rect 64880 9454 64932 9460
rect 64972 9512 65024 9518
rect 64972 9454 65024 9460
rect 64696 9172 64748 9178
rect 64696 9114 64748 9120
rect 64248 9030 64736 9058
rect 64236 8968 64288 8974
rect 64236 8910 64288 8916
rect 64052 7948 64104 7954
rect 64052 7890 64104 7896
rect 63960 6248 64012 6254
rect 63960 6190 64012 6196
rect 63960 5568 64012 5574
rect 63960 5510 64012 5516
rect 63868 4684 63920 4690
rect 63868 4626 63920 4632
rect 63972 4282 64000 5510
rect 64064 5234 64092 7890
rect 64142 6896 64198 6905
rect 64142 6831 64198 6840
rect 64156 6390 64184 6831
rect 64144 6384 64196 6390
rect 64144 6326 64196 6332
rect 64144 5908 64196 5914
rect 64144 5850 64196 5856
rect 64052 5228 64104 5234
rect 64052 5170 64104 5176
rect 63960 4276 64012 4282
rect 63960 4218 64012 4224
rect 64064 4010 64092 5170
rect 64156 4026 64184 5850
rect 64248 5794 64276 8910
rect 64338 8732 64646 8741
rect 64338 8730 64344 8732
rect 64400 8730 64424 8732
rect 64480 8730 64504 8732
rect 64560 8730 64584 8732
rect 64640 8730 64646 8732
rect 64400 8678 64402 8730
rect 64582 8678 64584 8730
rect 64338 8676 64344 8678
rect 64400 8676 64424 8678
rect 64480 8676 64504 8678
rect 64560 8676 64584 8678
rect 64640 8676 64646 8678
rect 64338 8667 64646 8676
rect 64604 8288 64656 8294
rect 64604 8230 64656 8236
rect 64616 8022 64644 8230
rect 64604 8016 64656 8022
rect 64604 7958 64656 7964
rect 64338 7644 64646 7653
rect 64338 7642 64344 7644
rect 64400 7642 64424 7644
rect 64480 7642 64504 7644
rect 64560 7642 64584 7644
rect 64640 7642 64646 7644
rect 64400 7590 64402 7642
rect 64582 7590 64584 7642
rect 64338 7588 64344 7590
rect 64400 7588 64424 7590
rect 64480 7588 64504 7590
rect 64560 7588 64584 7590
rect 64640 7588 64646 7590
rect 64338 7579 64646 7588
rect 64510 7440 64566 7449
rect 64510 7375 64566 7384
rect 64524 7342 64552 7375
rect 64512 7336 64564 7342
rect 64512 7278 64564 7284
rect 64524 6866 64552 7278
rect 64602 6896 64658 6905
rect 64512 6860 64564 6866
rect 64602 6831 64604 6840
rect 64512 6802 64564 6808
rect 64656 6831 64658 6840
rect 64604 6802 64656 6808
rect 64338 6556 64646 6565
rect 64338 6554 64344 6556
rect 64400 6554 64424 6556
rect 64480 6554 64504 6556
rect 64560 6554 64584 6556
rect 64640 6554 64646 6556
rect 64400 6502 64402 6554
rect 64582 6502 64584 6554
rect 64338 6500 64344 6502
rect 64400 6500 64424 6502
rect 64480 6500 64504 6502
rect 64560 6500 64584 6502
rect 64640 6500 64646 6502
rect 64338 6491 64646 6500
rect 64512 6384 64564 6390
rect 64512 6326 64564 6332
rect 64524 6254 64552 6326
rect 64512 6248 64564 6254
rect 64512 6190 64564 6196
rect 64328 6112 64380 6118
rect 64328 6054 64380 6060
rect 64340 5914 64368 6054
rect 64524 5914 64552 6190
rect 64328 5908 64380 5914
rect 64328 5850 64380 5856
rect 64512 5908 64564 5914
rect 64512 5850 64564 5856
rect 64248 5766 64368 5794
rect 64340 5710 64368 5766
rect 64328 5704 64380 5710
rect 64328 5646 64380 5652
rect 64338 5468 64646 5477
rect 64338 5466 64344 5468
rect 64400 5466 64424 5468
rect 64480 5466 64504 5468
rect 64560 5466 64584 5468
rect 64640 5466 64646 5468
rect 64400 5414 64402 5466
rect 64582 5414 64584 5466
rect 64338 5412 64344 5414
rect 64400 5412 64424 5414
rect 64480 5412 64504 5414
rect 64560 5412 64584 5414
rect 64640 5412 64646 5414
rect 64338 5403 64646 5412
rect 64708 4978 64736 9030
rect 64892 7478 64920 9454
rect 65064 9444 65116 9450
rect 65064 9386 65116 9392
rect 64972 9376 65024 9382
rect 64972 9318 65024 9324
rect 64984 9042 65012 9318
rect 65076 9178 65104 9386
rect 65156 9376 65208 9382
rect 65156 9318 65208 9324
rect 65064 9172 65116 9178
rect 65064 9114 65116 9120
rect 64972 9036 65024 9042
rect 64972 8978 65024 8984
rect 65064 8968 65116 8974
rect 65064 8910 65116 8916
rect 65076 7546 65104 8910
rect 65064 7540 65116 7546
rect 65064 7482 65116 7488
rect 64880 7472 64932 7478
rect 64880 7414 64932 7420
rect 64892 6914 64920 7414
rect 64892 6886 65012 6914
rect 64984 6798 65012 6886
rect 65168 6866 65196 9318
rect 65258 9276 65566 9285
rect 65258 9274 65264 9276
rect 65320 9274 65344 9276
rect 65400 9274 65424 9276
rect 65480 9274 65504 9276
rect 65560 9274 65566 9276
rect 65320 9222 65322 9274
rect 65502 9222 65504 9274
rect 65258 9220 65264 9222
rect 65320 9220 65344 9222
rect 65400 9220 65424 9222
rect 65480 9220 65504 9222
rect 65560 9220 65566 9222
rect 65258 9211 65566 9220
rect 65248 8968 65300 8974
rect 65248 8910 65300 8916
rect 65260 8498 65288 8910
rect 65248 8492 65300 8498
rect 65248 8434 65300 8440
rect 65628 8430 65656 10678
rect 65720 8974 65748 10798
rect 65812 10606 65840 16186
rect 65904 15638 65932 19246
rect 65984 18760 66036 18766
rect 65984 18702 66036 18708
rect 65996 18086 66024 18702
rect 66088 18426 66116 36314
rect 66180 31929 66208 36790
rect 66260 34672 66312 34678
rect 66260 34614 66312 34620
rect 66166 31920 66222 31929
rect 66166 31855 66222 31864
rect 66168 31816 66220 31822
rect 66168 31758 66220 31764
rect 66180 20330 66208 31758
rect 66272 22234 66300 34614
rect 66364 33046 66392 43794
rect 66444 41200 66496 41206
rect 66444 41142 66496 41148
rect 66352 33040 66404 33046
rect 66352 32982 66404 32988
rect 66364 31754 66392 32982
rect 66456 31890 66484 41142
rect 66536 36780 66588 36786
rect 66536 36722 66588 36728
rect 66548 33590 66576 36722
rect 66536 33584 66588 33590
rect 66536 33526 66588 33532
rect 66444 31884 66496 31890
rect 66444 31826 66496 31832
rect 66364 31726 66484 31754
rect 66456 30122 66484 31726
rect 66444 30116 66496 30122
rect 66444 30058 66496 30064
rect 66456 29034 66484 30058
rect 66548 29646 66576 33526
rect 66536 29640 66588 29646
rect 66536 29582 66588 29588
rect 66444 29028 66496 29034
rect 66444 28970 66496 28976
rect 66548 26382 66576 29582
rect 66536 26376 66588 26382
rect 66536 26318 66588 26324
rect 66260 22228 66312 22234
rect 66260 22170 66312 22176
rect 66272 21486 66300 22170
rect 66260 21480 66312 21486
rect 66260 21422 66312 21428
rect 66168 20324 66220 20330
rect 66168 20266 66220 20272
rect 66168 19984 66220 19990
rect 66168 19926 66220 19932
rect 66076 18420 66128 18426
rect 66076 18362 66128 18368
rect 66180 18154 66208 19926
rect 66168 18148 66220 18154
rect 66168 18090 66220 18096
rect 65984 18080 66036 18086
rect 65984 18022 66036 18028
rect 65984 17740 66036 17746
rect 65984 17682 66036 17688
rect 65892 15632 65944 15638
rect 65892 15574 65944 15580
rect 65996 12442 66024 17682
rect 66076 16720 66128 16726
rect 66076 16662 66128 16668
rect 66088 12850 66116 16662
rect 66180 15978 66208 18090
rect 66168 15972 66220 15978
rect 66168 15914 66220 15920
rect 66076 12844 66128 12850
rect 66076 12786 66128 12792
rect 65984 12436 66036 12442
rect 65984 12378 66036 12384
rect 65892 11552 65944 11558
rect 65892 11494 65944 11500
rect 65800 10600 65852 10606
rect 65800 10542 65852 10548
rect 65708 8968 65760 8974
rect 65708 8910 65760 8916
rect 65616 8424 65668 8430
rect 65616 8366 65668 8372
rect 65258 8188 65566 8197
rect 65258 8186 65264 8188
rect 65320 8186 65344 8188
rect 65400 8186 65424 8188
rect 65480 8186 65504 8188
rect 65560 8186 65566 8188
rect 65320 8134 65322 8186
rect 65502 8134 65504 8186
rect 65258 8132 65264 8134
rect 65320 8132 65344 8134
rect 65400 8132 65424 8134
rect 65480 8132 65504 8134
rect 65560 8132 65566 8134
rect 65258 8123 65566 8132
rect 65616 7200 65668 7206
rect 65616 7142 65668 7148
rect 65258 7100 65566 7109
rect 65258 7098 65264 7100
rect 65320 7098 65344 7100
rect 65400 7098 65424 7100
rect 65480 7098 65504 7100
rect 65560 7098 65566 7100
rect 65320 7046 65322 7098
rect 65502 7046 65504 7098
rect 65258 7044 65264 7046
rect 65320 7044 65344 7046
rect 65400 7044 65424 7046
rect 65480 7044 65504 7046
rect 65560 7044 65566 7046
rect 65258 7035 65566 7044
rect 65628 7002 65656 7142
rect 65616 6996 65668 7002
rect 65616 6938 65668 6944
rect 65156 6860 65208 6866
rect 65156 6802 65208 6808
rect 64972 6792 65024 6798
rect 64972 6734 65024 6740
rect 65616 6792 65668 6798
rect 65720 6746 65748 8910
rect 65800 8424 65852 8430
rect 65800 8366 65852 8372
rect 65812 7750 65840 8366
rect 65800 7744 65852 7750
rect 65800 7686 65852 7692
rect 65812 7410 65840 7686
rect 65800 7404 65852 7410
rect 65800 7346 65852 7352
rect 65668 6740 65748 6746
rect 65616 6734 65748 6740
rect 64788 6656 64840 6662
rect 64788 6598 64840 6604
rect 64800 5234 64828 6598
rect 64984 6322 65012 6734
rect 65628 6718 65748 6734
rect 64972 6316 65024 6322
rect 64972 6258 65024 6264
rect 64880 6180 64932 6186
rect 64880 6122 64932 6128
rect 64788 5228 64840 5234
rect 64788 5170 64840 5176
rect 64708 4950 64828 4978
rect 64696 4616 64748 4622
rect 64696 4558 64748 4564
rect 64338 4380 64646 4389
rect 64338 4378 64344 4380
rect 64400 4378 64424 4380
rect 64480 4378 64504 4380
rect 64560 4378 64584 4380
rect 64640 4378 64646 4380
rect 64400 4326 64402 4378
rect 64582 4326 64584 4378
rect 64338 4324 64344 4326
rect 64400 4324 64424 4326
rect 64480 4324 64504 4326
rect 64560 4324 64584 4326
rect 64640 4324 64646 4326
rect 64338 4315 64646 4324
rect 64052 4004 64104 4010
rect 64156 3998 64276 4026
rect 64052 3946 64104 3952
rect 63868 3664 63920 3670
rect 63868 3606 63920 3612
rect 63880 3194 63908 3606
rect 63868 3188 63920 3194
rect 63868 3130 63920 3136
rect 64064 3058 64092 3946
rect 64144 3936 64196 3942
rect 64144 3878 64196 3884
rect 64156 3738 64184 3878
rect 64144 3732 64196 3738
rect 64144 3674 64196 3680
rect 64052 3052 64104 3058
rect 64052 2994 64104 3000
rect 64156 2514 64184 3674
rect 64248 3074 64276 3998
rect 64708 3398 64736 4558
rect 64696 3392 64748 3398
rect 64696 3334 64748 3340
rect 64338 3292 64646 3301
rect 64338 3290 64344 3292
rect 64400 3290 64424 3292
rect 64480 3290 64504 3292
rect 64560 3290 64584 3292
rect 64640 3290 64646 3292
rect 64400 3238 64402 3290
rect 64582 3238 64584 3290
rect 64338 3236 64344 3238
rect 64400 3236 64424 3238
rect 64480 3236 64504 3238
rect 64560 3236 64584 3238
rect 64640 3236 64646 3238
rect 64338 3227 64646 3236
rect 64800 3074 64828 4950
rect 64892 4826 64920 6122
rect 64880 4820 64932 4826
rect 64880 4762 64932 4768
rect 64984 3466 65012 6258
rect 65258 6012 65566 6021
rect 65258 6010 65264 6012
rect 65320 6010 65344 6012
rect 65400 6010 65424 6012
rect 65480 6010 65504 6012
rect 65560 6010 65566 6012
rect 65320 5958 65322 6010
rect 65502 5958 65504 6010
rect 65258 5956 65264 5958
rect 65320 5956 65344 5958
rect 65400 5956 65424 5958
rect 65480 5956 65504 5958
rect 65560 5956 65566 5958
rect 65258 5947 65566 5956
rect 65258 4924 65566 4933
rect 65258 4922 65264 4924
rect 65320 4922 65344 4924
rect 65400 4922 65424 4924
rect 65480 4922 65504 4924
rect 65560 4922 65566 4924
rect 65320 4870 65322 4922
rect 65502 4870 65504 4922
rect 65258 4868 65264 4870
rect 65320 4868 65344 4870
rect 65400 4868 65424 4870
rect 65480 4868 65504 4870
rect 65560 4868 65566 4870
rect 65258 4859 65566 4868
rect 65156 4820 65208 4826
rect 65156 4762 65208 4768
rect 65064 3596 65116 3602
rect 65064 3538 65116 3544
rect 64972 3460 65024 3466
rect 64972 3402 65024 3408
rect 64248 3046 64368 3074
rect 64800 3046 65012 3074
rect 64236 2916 64288 2922
rect 64236 2858 64288 2864
rect 64144 2508 64196 2514
rect 64144 2450 64196 2456
rect 63776 1896 63828 1902
rect 63682 1864 63738 1873
rect 63776 1838 63828 1844
rect 63682 1799 63738 1808
rect 64248 1426 64276 2858
rect 64340 2446 64368 3046
rect 64984 2650 65012 3046
rect 64972 2644 65024 2650
rect 64972 2586 65024 2592
rect 64328 2440 64380 2446
rect 64328 2382 64380 2388
rect 64696 2440 64748 2446
rect 64696 2382 64748 2388
rect 64338 2204 64646 2213
rect 64338 2202 64344 2204
rect 64400 2202 64424 2204
rect 64480 2202 64504 2204
rect 64560 2202 64584 2204
rect 64640 2202 64646 2204
rect 64400 2150 64402 2202
rect 64582 2150 64584 2202
rect 64338 2148 64344 2150
rect 64400 2148 64424 2150
rect 64480 2148 64504 2150
rect 64560 2148 64584 2150
rect 64640 2148 64646 2150
rect 64338 2139 64646 2148
rect 64708 1970 64736 2382
rect 64788 2304 64840 2310
rect 64788 2246 64840 2252
rect 64696 1964 64748 1970
rect 64696 1906 64748 1912
rect 64696 1828 64748 1834
rect 64696 1770 64748 1776
rect 64708 1562 64736 1770
rect 64800 1562 64828 2246
rect 64984 1834 65012 2586
rect 65076 2106 65104 3538
rect 65168 2514 65196 4762
rect 65258 3836 65566 3845
rect 65258 3834 65264 3836
rect 65320 3834 65344 3836
rect 65400 3834 65424 3836
rect 65480 3834 65504 3836
rect 65560 3834 65566 3836
rect 65320 3782 65322 3834
rect 65502 3782 65504 3834
rect 65258 3780 65264 3782
rect 65320 3780 65344 3782
rect 65400 3780 65424 3782
rect 65480 3780 65504 3782
rect 65560 3780 65566 3782
rect 65258 3771 65566 3780
rect 65628 3534 65656 6718
rect 65708 5092 65760 5098
rect 65708 5034 65760 5040
rect 65720 4758 65748 5034
rect 65708 4752 65760 4758
rect 65708 4694 65760 4700
rect 65616 3528 65668 3534
rect 65616 3470 65668 3476
rect 65258 2748 65566 2757
rect 65258 2746 65264 2748
rect 65320 2746 65344 2748
rect 65400 2746 65424 2748
rect 65480 2746 65504 2748
rect 65560 2746 65566 2748
rect 65320 2694 65322 2746
rect 65502 2694 65504 2746
rect 65258 2692 65264 2694
rect 65320 2692 65344 2694
rect 65400 2692 65424 2694
rect 65480 2692 65504 2694
rect 65560 2692 65566 2694
rect 65258 2683 65566 2692
rect 65156 2508 65208 2514
rect 65156 2450 65208 2456
rect 65064 2100 65116 2106
rect 65064 2042 65116 2048
rect 65168 1902 65196 2450
rect 65156 1896 65208 1902
rect 65156 1838 65208 1844
rect 64972 1828 65024 1834
rect 64972 1770 65024 1776
rect 65258 1660 65566 1669
rect 65258 1658 65264 1660
rect 65320 1658 65344 1660
rect 65400 1658 65424 1660
rect 65480 1658 65504 1660
rect 65560 1658 65566 1660
rect 65320 1606 65322 1658
rect 65502 1606 65504 1658
rect 65258 1604 65264 1606
rect 65320 1604 65344 1606
rect 65400 1604 65424 1606
rect 65480 1604 65504 1606
rect 65560 1604 65566 1606
rect 65258 1595 65566 1604
rect 64696 1556 64748 1562
rect 64696 1498 64748 1504
rect 64788 1556 64840 1562
rect 64788 1498 64840 1504
rect 64236 1420 64288 1426
rect 64236 1362 64288 1368
rect 65156 1420 65208 1426
rect 65156 1362 65208 1368
rect 62946 1320 63002 1329
rect 62946 1255 63002 1264
rect 64338 1116 64646 1125
rect 64338 1114 64344 1116
rect 64400 1114 64424 1116
rect 64480 1114 64504 1116
rect 64560 1114 64584 1116
rect 64640 1114 64646 1116
rect 64400 1062 64402 1114
rect 64582 1062 64584 1114
rect 64338 1060 64344 1062
rect 64400 1060 64424 1062
rect 64480 1060 64504 1062
rect 64560 1060 64584 1062
rect 64640 1060 64646 1062
rect 64338 1051 64646 1060
rect 65168 1018 65196 1362
rect 65628 1358 65656 3470
rect 65720 2922 65748 4694
rect 65708 2916 65760 2922
rect 65708 2858 65760 2864
rect 65800 2848 65852 2854
rect 65800 2790 65852 2796
rect 65812 1970 65840 2790
rect 65904 2038 65932 11494
rect 65996 11218 66024 12378
rect 66088 11626 66116 12786
rect 66180 12374 66208 15914
rect 66444 12640 66496 12646
rect 66444 12582 66496 12588
rect 66168 12368 66220 12374
rect 66168 12310 66220 12316
rect 66076 11620 66128 11626
rect 66076 11562 66128 11568
rect 65984 11212 66036 11218
rect 65984 11154 66036 11160
rect 65996 9042 66024 11154
rect 65984 9036 66036 9042
rect 65984 8978 66036 8984
rect 65984 7336 66036 7342
rect 65984 7278 66036 7284
rect 65996 6254 66024 7278
rect 65984 6248 66036 6254
rect 65984 6190 66036 6196
rect 65996 5370 66024 6190
rect 65984 5364 66036 5370
rect 65984 5306 66036 5312
rect 66088 2650 66116 11562
rect 66180 10198 66208 12310
rect 66260 11688 66312 11694
rect 66260 11630 66312 11636
rect 66168 10192 66220 10198
rect 66168 10134 66220 10140
rect 66180 8022 66208 10134
rect 66168 8016 66220 8022
rect 66168 7958 66220 7964
rect 66180 5098 66208 7958
rect 66272 6458 66300 11630
rect 66260 6452 66312 6458
rect 66260 6394 66312 6400
rect 66168 5092 66220 5098
rect 66168 5034 66220 5040
rect 66456 4010 66484 12582
rect 66444 4004 66496 4010
rect 66444 3946 66496 3952
rect 66076 2644 66128 2650
rect 66076 2586 66128 2592
rect 65892 2032 65944 2038
rect 65892 1974 65944 1980
rect 65800 1964 65852 1970
rect 65800 1906 65852 1912
rect 65616 1352 65668 1358
rect 65616 1294 65668 1300
rect 65156 1012 65208 1018
rect 65156 954 65208 960
rect 65812 882 65840 1906
rect 65800 876 65852 882
rect 65800 818 65852 824
rect 65258 572 65566 581
rect 65258 570 65264 572
rect 65320 570 65344 572
rect 65400 570 65424 572
rect 65480 570 65504 572
rect 65560 570 65566 572
rect 65320 518 65322 570
rect 65502 518 65504 570
rect 65258 516 65264 518
rect 65320 516 65344 518
rect 65400 516 65424 518
rect 65480 516 65504 518
rect 65560 516 65566 518
rect 65258 507 65566 516
<< via2 >>
rect 34610 45056 34666 45112
rect 11702 44784 11758 44840
rect 13818 44784 13874 44840
rect 11150 44648 11206 44704
rect 2004 44634 2060 44636
rect 2084 44634 2140 44636
rect 2164 44634 2220 44636
rect 2244 44634 2300 44636
rect 2004 44582 2050 44634
rect 2050 44582 2060 44634
rect 2084 44582 2114 44634
rect 2114 44582 2126 44634
rect 2126 44582 2140 44634
rect 2164 44582 2178 44634
rect 2178 44582 2190 44634
rect 2190 44582 2220 44634
rect 2244 44582 2254 44634
rect 2254 44582 2300 44634
rect 2004 44580 2060 44582
rect 2084 44580 2140 44582
rect 2164 44580 2220 44582
rect 2244 44580 2300 44582
rect 6182 44532 6238 44568
rect 6182 44512 6184 44532
rect 6184 44512 6236 44532
rect 6236 44512 6238 44532
rect 6734 44532 6790 44568
rect 6734 44512 6736 44532
rect 6736 44512 6788 44532
rect 6788 44512 6790 44532
rect 7286 44532 7342 44568
rect 7286 44512 7288 44532
rect 7288 44512 7340 44532
rect 7340 44512 7342 44532
rect 7838 44532 7894 44568
rect 7838 44512 7840 44532
rect 7840 44512 7892 44532
rect 7892 44512 7894 44532
rect 8390 44532 8446 44568
rect 8390 44512 8392 44532
rect 8392 44512 8444 44532
rect 8444 44512 8446 44532
rect 8942 44532 8998 44568
rect 8942 44512 8944 44532
rect 8944 44512 8996 44532
rect 8996 44512 8998 44532
rect 9494 44532 9550 44568
rect 9494 44512 9496 44532
rect 9496 44512 9548 44532
rect 9548 44512 9550 44532
rect 10046 44532 10102 44568
rect 10046 44512 10048 44532
rect 10048 44512 10100 44532
rect 10100 44512 10102 44532
rect 10506 44532 10562 44568
rect 10506 44512 10508 44532
rect 10508 44512 10560 44532
rect 10560 44512 10562 44532
rect 10782 44532 10838 44568
rect 10782 44512 10784 44532
rect 10784 44512 10836 44532
rect 10836 44512 10838 44532
rect 11426 44532 11482 44568
rect 11426 44512 11428 44532
rect 11428 44512 11480 44532
rect 11480 44512 11482 44532
rect 12530 44532 12586 44568
rect 12530 44512 12532 44532
rect 12532 44512 12584 44532
rect 12584 44512 12586 44532
rect 14370 44648 14426 44704
rect 15198 44532 15254 44568
rect 15198 44512 15200 44532
rect 15200 44512 15252 44532
rect 15252 44512 15254 44532
rect 20074 44532 20130 44568
rect 20074 44512 20076 44532
rect 20076 44512 20128 44532
rect 20128 44512 20130 44532
rect 2924 44090 2980 44092
rect 3004 44090 3060 44092
rect 3084 44090 3140 44092
rect 3164 44090 3220 44092
rect 2924 44038 2970 44090
rect 2970 44038 2980 44090
rect 3004 44038 3034 44090
rect 3034 44038 3046 44090
rect 3046 44038 3060 44090
rect 3084 44038 3098 44090
rect 3098 44038 3110 44090
rect 3110 44038 3140 44090
rect 3164 44038 3174 44090
rect 3174 44038 3220 44090
rect 2924 44036 2980 44038
rect 3004 44036 3060 44038
rect 3084 44036 3140 44038
rect 3164 44036 3220 44038
rect 2004 43546 2060 43548
rect 2084 43546 2140 43548
rect 2164 43546 2220 43548
rect 2244 43546 2300 43548
rect 2004 43494 2050 43546
rect 2050 43494 2060 43546
rect 2084 43494 2114 43546
rect 2114 43494 2126 43546
rect 2126 43494 2140 43546
rect 2164 43494 2178 43546
rect 2178 43494 2190 43546
rect 2190 43494 2220 43546
rect 2244 43494 2254 43546
rect 2254 43494 2300 43546
rect 2004 43492 2060 43494
rect 2084 43492 2140 43494
rect 2164 43492 2220 43494
rect 2244 43492 2300 43494
rect 2924 43002 2980 43004
rect 3004 43002 3060 43004
rect 3084 43002 3140 43004
rect 3164 43002 3220 43004
rect 2924 42950 2970 43002
rect 2970 42950 2980 43002
rect 3004 42950 3034 43002
rect 3034 42950 3046 43002
rect 3046 42950 3060 43002
rect 3084 42950 3098 43002
rect 3098 42950 3110 43002
rect 3110 42950 3140 43002
rect 3164 42950 3174 43002
rect 3174 42950 3220 43002
rect 2924 42948 2980 42950
rect 3004 42948 3060 42950
rect 3084 42948 3140 42950
rect 3164 42948 3220 42950
rect 2004 42458 2060 42460
rect 2084 42458 2140 42460
rect 2164 42458 2220 42460
rect 2244 42458 2300 42460
rect 2004 42406 2050 42458
rect 2050 42406 2060 42458
rect 2084 42406 2114 42458
rect 2114 42406 2126 42458
rect 2126 42406 2140 42458
rect 2164 42406 2178 42458
rect 2178 42406 2190 42458
rect 2190 42406 2220 42458
rect 2244 42406 2254 42458
rect 2254 42406 2300 42458
rect 2004 42404 2060 42406
rect 2084 42404 2140 42406
rect 2164 42404 2220 42406
rect 2244 42404 2300 42406
rect 2924 41914 2980 41916
rect 3004 41914 3060 41916
rect 3084 41914 3140 41916
rect 3164 41914 3220 41916
rect 2924 41862 2970 41914
rect 2970 41862 2980 41914
rect 3004 41862 3034 41914
rect 3034 41862 3046 41914
rect 3046 41862 3060 41914
rect 3084 41862 3098 41914
rect 3098 41862 3110 41914
rect 3110 41862 3140 41914
rect 3164 41862 3174 41914
rect 3174 41862 3220 41914
rect 2924 41860 2980 41862
rect 3004 41860 3060 41862
rect 3084 41860 3140 41862
rect 3164 41860 3220 41862
rect 2004 41370 2060 41372
rect 2084 41370 2140 41372
rect 2164 41370 2220 41372
rect 2244 41370 2300 41372
rect 2004 41318 2050 41370
rect 2050 41318 2060 41370
rect 2084 41318 2114 41370
rect 2114 41318 2126 41370
rect 2126 41318 2140 41370
rect 2164 41318 2178 41370
rect 2178 41318 2190 41370
rect 2190 41318 2220 41370
rect 2244 41318 2254 41370
rect 2254 41318 2300 41370
rect 2004 41316 2060 41318
rect 2084 41316 2140 41318
rect 2164 41316 2220 41318
rect 2244 41316 2300 41318
rect 2924 40826 2980 40828
rect 3004 40826 3060 40828
rect 3084 40826 3140 40828
rect 3164 40826 3220 40828
rect 2924 40774 2970 40826
rect 2970 40774 2980 40826
rect 3004 40774 3034 40826
rect 3034 40774 3046 40826
rect 3046 40774 3060 40826
rect 3084 40774 3098 40826
rect 3098 40774 3110 40826
rect 3110 40774 3140 40826
rect 3164 40774 3174 40826
rect 3174 40774 3220 40826
rect 2924 40772 2980 40774
rect 3004 40772 3060 40774
rect 3084 40772 3140 40774
rect 3164 40772 3220 40774
rect 2004 40282 2060 40284
rect 2084 40282 2140 40284
rect 2164 40282 2220 40284
rect 2244 40282 2300 40284
rect 2004 40230 2050 40282
rect 2050 40230 2060 40282
rect 2084 40230 2114 40282
rect 2114 40230 2126 40282
rect 2126 40230 2140 40282
rect 2164 40230 2178 40282
rect 2178 40230 2190 40282
rect 2190 40230 2220 40282
rect 2244 40230 2254 40282
rect 2254 40230 2300 40282
rect 2004 40228 2060 40230
rect 2084 40228 2140 40230
rect 2164 40228 2220 40230
rect 2244 40228 2300 40230
rect 2924 39738 2980 39740
rect 3004 39738 3060 39740
rect 3084 39738 3140 39740
rect 3164 39738 3220 39740
rect 2924 39686 2970 39738
rect 2970 39686 2980 39738
rect 3004 39686 3034 39738
rect 3034 39686 3046 39738
rect 3046 39686 3060 39738
rect 3084 39686 3098 39738
rect 3098 39686 3110 39738
rect 3110 39686 3140 39738
rect 3164 39686 3174 39738
rect 3174 39686 3220 39738
rect 2924 39684 2980 39686
rect 3004 39684 3060 39686
rect 3084 39684 3140 39686
rect 3164 39684 3220 39686
rect 2004 39194 2060 39196
rect 2084 39194 2140 39196
rect 2164 39194 2220 39196
rect 2244 39194 2300 39196
rect 2004 39142 2050 39194
rect 2050 39142 2060 39194
rect 2084 39142 2114 39194
rect 2114 39142 2126 39194
rect 2126 39142 2140 39194
rect 2164 39142 2178 39194
rect 2178 39142 2190 39194
rect 2190 39142 2220 39194
rect 2244 39142 2254 39194
rect 2254 39142 2300 39194
rect 2004 39140 2060 39142
rect 2084 39140 2140 39142
rect 2164 39140 2220 39142
rect 2244 39140 2300 39142
rect 2924 38650 2980 38652
rect 3004 38650 3060 38652
rect 3084 38650 3140 38652
rect 3164 38650 3220 38652
rect 2924 38598 2970 38650
rect 2970 38598 2980 38650
rect 3004 38598 3034 38650
rect 3034 38598 3046 38650
rect 3046 38598 3060 38650
rect 3084 38598 3098 38650
rect 3098 38598 3110 38650
rect 3110 38598 3140 38650
rect 3164 38598 3174 38650
rect 3174 38598 3220 38650
rect 2924 38596 2980 38598
rect 3004 38596 3060 38598
rect 3084 38596 3140 38598
rect 3164 38596 3220 38598
rect 2004 38106 2060 38108
rect 2084 38106 2140 38108
rect 2164 38106 2220 38108
rect 2244 38106 2300 38108
rect 2004 38054 2050 38106
rect 2050 38054 2060 38106
rect 2084 38054 2114 38106
rect 2114 38054 2126 38106
rect 2126 38054 2140 38106
rect 2164 38054 2178 38106
rect 2178 38054 2190 38106
rect 2190 38054 2220 38106
rect 2244 38054 2254 38106
rect 2254 38054 2300 38106
rect 2004 38052 2060 38054
rect 2084 38052 2140 38054
rect 2164 38052 2220 38054
rect 2244 38052 2300 38054
rect 2924 37562 2980 37564
rect 3004 37562 3060 37564
rect 3084 37562 3140 37564
rect 3164 37562 3220 37564
rect 2924 37510 2970 37562
rect 2970 37510 2980 37562
rect 3004 37510 3034 37562
rect 3034 37510 3046 37562
rect 3046 37510 3060 37562
rect 3084 37510 3098 37562
rect 3098 37510 3110 37562
rect 3110 37510 3140 37562
rect 3164 37510 3174 37562
rect 3174 37510 3220 37562
rect 2924 37508 2980 37510
rect 3004 37508 3060 37510
rect 3084 37508 3140 37510
rect 3164 37508 3220 37510
rect 11426 39616 11482 39672
rect 12806 43852 12862 43888
rect 12806 43832 12808 43852
rect 12808 43832 12860 43852
rect 12860 43832 12862 43852
rect 2004 37018 2060 37020
rect 2084 37018 2140 37020
rect 2164 37018 2220 37020
rect 2244 37018 2300 37020
rect 2004 36966 2050 37018
rect 2050 36966 2060 37018
rect 2084 36966 2114 37018
rect 2114 36966 2126 37018
rect 2126 36966 2140 37018
rect 2164 36966 2178 37018
rect 2178 36966 2190 37018
rect 2190 36966 2220 37018
rect 2244 36966 2254 37018
rect 2254 36966 2300 37018
rect 2004 36964 2060 36966
rect 2084 36964 2140 36966
rect 2164 36964 2220 36966
rect 2244 36964 2300 36966
rect 14002 40996 14058 41032
rect 14002 40976 14004 40996
rect 14004 40976 14056 40996
rect 14056 40976 14058 40996
rect 13634 39888 13690 39944
rect 12622 37440 12678 37496
rect 16210 43852 16266 43888
rect 16210 43832 16212 43852
rect 16212 43832 16264 43852
rect 16264 43832 16266 43852
rect 15566 42200 15622 42256
rect 17498 43444 17554 43480
rect 17498 43424 17500 43444
rect 17500 43424 17552 43444
rect 17552 43424 17554 43444
rect 17314 42880 17370 42936
rect 17958 42336 18014 42392
rect 16210 38800 16266 38856
rect 16210 36896 16266 36952
rect 18326 43988 18382 44024
rect 18326 43968 18328 43988
rect 18328 43968 18380 43988
rect 18380 43968 18382 43988
rect 17958 42084 18014 42120
rect 17958 42064 17960 42084
rect 17960 42064 18012 42084
rect 18012 42064 18014 42084
rect 20442 43152 20498 43208
rect 16578 37848 16634 37904
rect 27986 44784 28042 44840
rect 21362 42644 21364 42664
rect 21364 42644 21416 42664
rect 21416 42644 21418 42664
rect 21362 42608 21418 42644
rect 18510 40296 18566 40352
rect 12346 36624 12402 36680
rect 16394 36624 16450 36680
rect 18050 37712 18106 37768
rect 17958 37576 18014 37632
rect 17958 36488 18014 36544
rect 17866 35944 17922 36000
rect 8206 35672 8262 35728
rect 8482 35672 8538 35728
rect 20810 40432 20866 40488
rect 22098 41656 22154 41712
rect 21178 39208 21234 39264
rect 21086 38936 21142 38992
rect 19338 36896 19394 36952
rect 20718 36760 20774 36816
rect 21086 37168 21142 37224
rect 21178 37032 21234 37088
rect 20994 35944 21050 36000
rect 20626 35808 20682 35864
rect 22374 41656 22430 41712
rect 27342 44648 27398 44704
rect 23110 41656 23166 41712
rect 22650 40840 22706 40896
rect 24214 42608 24270 42664
rect 25686 44396 25742 44432
rect 25686 44376 25688 44396
rect 25688 44376 25740 44396
rect 25740 44376 25742 44396
rect 24950 43016 25006 43072
rect 25318 42608 25374 42664
rect 25226 41928 25282 41984
rect 24674 41520 24730 41576
rect 25042 40024 25098 40080
rect 25042 39480 25098 39536
rect 25042 39208 25098 39264
rect 24582 38548 24638 38584
rect 24582 38528 24584 38548
rect 24584 38528 24636 38548
rect 24636 38528 24638 38548
rect 23478 37168 23534 37224
rect 23202 36760 23258 36816
rect 25502 43016 25558 43072
rect 25962 43560 26018 43616
rect 25502 41792 25558 41848
rect 25410 36080 25466 36136
rect 24674 35980 24676 36000
rect 24676 35980 24728 36000
rect 24728 35980 24730 36000
rect 24674 35944 24730 35980
rect 23202 35808 23258 35864
rect 26146 42880 26202 42936
rect 28722 44648 28778 44704
rect 25778 41656 25834 41712
rect 26054 41656 26110 41712
rect 25870 41248 25926 41304
rect 26054 41384 26110 41440
rect 25962 40976 26018 41032
rect 26146 40976 26202 41032
rect 25778 37440 25834 37496
rect 26606 38664 26662 38720
rect 26698 38120 26754 38176
rect 26698 37712 26754 37768
rect 27618 39616 27674 39672
rect 27434 38528 27490 38584
rect 27526 37576 27582 37632
rect 27802 37848 27858 37904
rect 27986 38936 28042 38992
rect 28538 38392 28594 38448
rect 28354 38120 28410 38176
rect 28078 37732 28134 37768
rect 28078 37712 28080 37732
rect 28080 37712 28132 37732
rect 28132 37712 28134 37732
rect 28354 37712 28410 37768
rect 28538 38120 28594 38176
rect 28354 37440 28410 37496
rect 28538 37440 28594 37496
rect 27526 36488 27582 36544
rect 27250 36352 27306 36408
rect 27618 36216 27674 36272
rect 29642 41928 29698 41984
rect 29182 41676 29238 41712
rect 29182 41656 29184 41676
rect 29184 41656 29236 41676
rect 29236 41656 29238 41676
rect 30378 41656 30434 41712
rect 30378 41520 30434 41576
rect 30378 41112 30434 41168
rect 30654 42064 30710 42120
rect 30654 41928 30710 41984
rect 30654 41248 30710 41304
rect 30378 39072 30434 39128
rect 28906 37460 28962 37496
rect 28906 37440 28908 37460
rect 28908 37440 28960 37460
rect 28960 37440 28962 37460
rect 28998 37304 29054 37360
rect 28630 37168 28686 37224
rect 20074 35672 20130 35728
rect 21178 35672 21234 35728
rect 22006 35672 22062 35728
rect 22190 35672 22246 35728
rect 25502 35808 25558 35864
rect 25870 35808 25926 35864
rect 30838 38528 30894 38584
rect 30838 37848 30894 37904
rect 30654 35944 30710 36000
rect 30930 35944 30986 36000
rect 23018 35708 23020 35728
rect 23020 35708 23072 35728
rect 23072 35708 23074 35728
rect 23018 35672 23074 35708
rect 23570 35672 23626 35728
rect 30286 35808 30342 35864
rect 31298 40160 31354 40216
rect 34242 43288 34298 43344
rect 32034 42064 32090 42120
rect 31390 38936 31446 38992
rect 31574 39208 31630 39264
rect 31482 37848 31538 37904
rect 31850 39888 31906 39944
rect 33322 41112 33378 41168
rect 34426 40568 34482 40624
rect 33046 38936 33102 38992
rect 31942 38664 31998 38720
rect 32126 38664 32182 38720
rect 32310 37460 32366 37496
rect 32310 37440 32312 37460
rect 32312 37440 32364 37460
rect 32364 37440 32366 37460
rect 33230 38412 33286 38448
rect 33230 38392 33232 38412
rect 33232 38392 33284 38412
rect 33284 38392 33286 38412
rect 33138 38120 33194 38176
rect 33230 37712 33286 37768
rect 33138 37440 33194 37496
rect 33598 38664 33654 38720
rect 33690 38120 33746 38176
rect 33690 37712 33746 37768
rect 33414 36080 33470 36136
rect 34426 39752 34482 39808
rect 34794 41384 34850 41440
rect 34702 40024 34758 40080
rect 36174 43016 36230 43072
rect 35898 42200 35954 42256
rect 34242 37868 34298 37904
rect 34242 37848 34244 37868
rect 34244 37848 34296 37868
rect 34296 37848 34298 37868
rect 34702 37712 34758 37768
rect 34978 38528 35034 38584
rect 35806 39888 35862 39944
rect 35622 38528 35678 38584
rect 35346 37576 35402 37632
rect 35438 37440 35494 37496
rect 37094 42336 37150 42392
rect 36726 40976 36782 41032
rect 36634 39616 36690 39672
rect 35530 36216 35586 36272
rect 31666 35808 31722 35864
rect 34150 35808 34206 35864
rect 34426 35808 34482 35864
rect 36726 39208 36782 39264
rect 50004 44634 50060 44636
rect 50084 44634 50140 44636
rect 50164 44634 50220 44636
rect 50244 44634 50300 44636
rect 50004 44582 50050 44634
rect 50050 44582 50060 44634
rect 50084 44582 50114 44634
rect 50114 44582 50126 44634
rect 50126 44582 50140 44634
rect 50164 44582 50178 44634
rect 50178 44582 50190 44634
rect 50190 44582 50220 44634
rect 50244 44582 50254 44634
rect 50254 44582 50300 44634
rect 50004 44580 50060 44582
rect 50084 44580 50140 44582
rect 50164 44580 50220 44582
rect 50244 44580 50300 44582
rect 37186 37168 37242 37224
rect 38842 40160 38898 40216
rect 38750 39616 38806 39672
rect 37738 36760 37794 36816
rect 36542 36488 36598 36544
rect 41786 43052 41788 43072
rect 41788 43052 41840 43072
rect 41840 43052 41842 43072
rect 41786 43016 41842 43052
rect 40682 41248 40738 41304
rect 39670 37848 39726 37904
rect 41050 39788 41052 39808
rect 41052 39788 41104 39808
rect 41104 39788 41106 39808
rect 41050 39752 41106 39788
rect 41970 40704 42026 40760
rect 43074 41792 43130 41848
rect 41234 39208 41290 39264
rect 41050 38528 41106 38584
rect 41326 37848 41382 37904
rect 41602 39208 41658 39264
rect 41970 38256 42026 38312
rect 39394 37032 39450 37088
rect 38658 36216 38714 36272
rect 38658 36100 38714 36136
rect 38658 36080 38660 36100
rect 38660 36080 38712 36100
rect 38712 36080 38714 36100
rect 35806 35964 35862 36000
rect 35806 35944 35808 35964
rect 35808 35944 35860 35964
rect 35860 35944 35862 35964
rect 44270 43016 44326 43072
rect 43534 41656 43590 41712
rect 44270 42084 44326 42120
rect 44270 42064 44272 42084
rect 44272 42064 44324 42084
rect 44324 42064 44326 42084
rect 43902 41248 43958 41304
rect 44730 39752 44786 39808
rect 43902 38664 43958 38720
rect 45098 39380 45100 39400
rect 45100 39380 45152 39400
rect 45152 39380 45154 39400
rect 45098 39344 45154 39380
rect 44546 38004 44602 38040
rect 44546 37984 44548 38004
rect 44548 37984 44600 38004
rect 44600 37984 44602 38004
rect 45098 38528 45154 38584
rect 47398 42608 47454 42664
rect 50924 44090 50980 44092
rect 51004 44090 51060 44092
rect 51084 44090 51140 44092
rect 51164 44090 51220 44092
rect 50924 44038 50970 44090
rect 50970 44038 50980 44090
rect 51004 44038 51034 44090
rect 51034 44038 51046 44090
rect 51046 44038 51060 44090
rect 51084 44038 51098 44090
rect 51098 44038 51110 44090
rect 51110 44038 51140 44090
rect 51164 44038 51174 44090
rect 51174 44038 51220 44090
rect 50924 44036 50980 44038
rect 51004 44036 51060 44038
rect 51084 44036 51140 44038
rect 51164 44036 51220 44038
rect 50004 43546 50060 43548
rect 50084 43546 50140 43548
rect 50164 43546 50220 43548
rect 50244 43546 50300 43548
rect 50004 43494 50050 43546
rect 50050 43494 50060 43546
rect 50084 43494 50114 43546
rect 50114 43494 50126 43546
rect 50126 43494 50140 43546
rect 50164 43494 50178 43546
rect 50178 43494 50190 43546
rect 50190 43494 50220 43546
rect 50244 43494 50254 43546
rect 50254 43494 50300 43546
rect 50004 43492 50060 43494
rect 50084 43492 50140 43494
rect 50164 43492 50220 43494
rect 50244 43492 50300 43494
rect 47858 40588 47914 40624
rect 47858 40568 47860 40588
rect 47860 40568 47912 40588
rect 47912 40568 47914 40588
rect 48226 40568 48282 40624
rect 48318 38528 48374 38584
rect 50924 43002 50980 43004
rect 51004 43002 51060 43004
rect 51084 43002 51140 43004
rect 51164 43002 51220 43004
rect 50924 42950 50970 43002
rect 50970 42950 50980 43002
rect 51004 42950 51034 43002
rect 51034 42950 51046 43002
rect 51046 42950 51060 43002
rect 51084 42950 51098 43002
rect 51098 42950 51110 43002
rect 51110 42950 51140 43002
rect 51164 42950 51174 43002
rect 51174 42950 51220 43002
rect 50924 42948 50980 42950
rect 51004 42948 51060 42950
rect 51084 42948 51140 42950
rect 51164 42948 51220 42950
rect 50004 42458 50060 42460
rect 50084 42458 50140 42460
rect 50164 42458 50220 42460
rect 50244 42458 50300 42460
rect 50004 42406 50050 42458
rect 50050 42406 50060 42458
rect 50084 42406 50114 42458
rect 50114 42406 50126 42458
rect 50126 42406 50140 42458
rect 50164 42406 50178 42458
rect 50178 42406 50190 42458
rect 50190 42406 50220 42458
rect 50244 42406 50254 42458
rect 50254 42406 50300 42458
rect 50004 42404 50060 42406
rect 50084 42404 50140 42406
rect 50164 42404 50220 42406
rect 50244 42404 50300 42406
rect 49790 40432 49846 40488
rect 50004 41370 50060 41372
rect 50084 41370 50140 41372
rect 50164 41370 50220 41372
rect 50244 41370 50300 41372
rect 50004 41318 50050 41370
rect 50050 41318 50060 41370
rect 50084 41318 50114 41370
rect 50114 41318 50126 41370
rect 50126 41318 50140 41370
rect 50164 41318 50178 41370
rect 50178 41318 50190 41370
rect 50190 41318 50220 41370
rect 50244 41318 50254 41370
rect 50254 41318 50300 41370
rect 50004 41316 50060 41318
rect 50084 41316 50140 41318
rect 50164 41316 50220 41318
rect 50244 41316 50300 41318
rect 50924 41914 50980 41916
rect 51004 41914 51060 41916
rect 51084 41914 51140 41916
rect 51164 41914 51220 41916
rect 50924 41862 50970 41914
rect 50970 41862 50980 41914
rect 51004 41862 51034 41914
rect 51034 41862 51046 41914
rect 51046 41862 51060 41914
rect 51084 41862 51098 41914
rect 51098 41862 51110 41914
rect 51110 41862 51140 41914
rect 51164 41862 51174 41914
rect 51174 41862 51220 41914
rect 50924 41860 50980 41862
rect 51004 41860 51060 41862
rect 51084 41860 51140 41862
rect 51164 41860 51220 41862
rect 50894 40976 50950 41032
rect 50924 40826 50980 40828
rect 51004 40826 51060 40828
rect 51084 40826 51140 40828
rect 51164 40826 51220 40828
rect 50924 40774 50970 40826
rect 50970 40774 50980 40826
rect 51004 40774 51034 40826
rect 51034 40774 51046 40826
rect 51046 40774 51060 40826
rect 51084 40774 51098 40826
rect 51098 40774 51110 40826
rect 51110 40774 51140 40826
rect 51164 40774 51174 40826
rect 51174 40774 51220 40826
rect 50924 40772 50980 40774
rect 51004 40772 51060 40774
rect 51084 40772 51140 40774
rect 51164 40772 51220 40774
rect 50004 40282 50060 40284
rect 50084 40282 50140 40284
rect 50164 40282 50220 40284
rect 50244 40282 50300 40284
rect 50004 40230 50050 40282
rect 50050 40230 50060 40282
rect 50084 40230 50114 40282
rect 50114 40230 50126 40282
rect 50126 40230 50140 40282
rect 50164 40230 50178 40282
rect 50178 40230 50190 40282
rect 50190 40230 50220 40282
rect 50244 40230 50254 40282
rect 50254 40230 50300 40282
rect 50004 40228 50060 40230
rect 50084 40228 50140 40230
rect 50164 40228 50220 40230
rect 50244 40228 50300 40230
rect 50924 39738 50980 39740
rect 51004 39738 51060 39740
rect 51084 39738 51140 39740
rect 51164 39738 51220 39740
rect 50924 39686 50970 39738
rect 50970 39686 50980 39738
rect 51004 39686 51034 39738
rect 51034 39686 51046 39738
rect 51046 39686 51060 39738
rect 51084 39686 51098 39738
rect 51098 39686 51110 39738
rect 51110 39686 51140 39738
rect 51164 39686 51174 39738
rect 51174 39686 51220 39738
rect 50924 39684 50980 39686
rect 51004 39684 51060 39686
rect 51084 39684 51140 39686
rect 51164 39684 51220 39686
rect 50004 39194 50060 39196
rect 50084 39194 50140 39196
rect 50164 39194 50220 39196
rect 50244 39194 50300 39196
rect 50004 39142 50050 39194
rect 50050 39142 50060 39194
rect 50084 39142 50114 39194
rect 50114 39142 50126 39194
rect 50126 39142 50140 39194
rect 50164 39142 50178 39194
rect 50178 39142 50190 39194
rect 50190 39142 50220 39194
rect 50244 39142 50254 39194
rect 50254 39142 50300 39194
rect 50004 39140 50060 39142
rect 50084 39140 50140 39142
rect 50164 39140 50220 39142
rect 50244 39140 50300 39142
rect 48870 38528 48926 38584
rect 48410 37304 48466 37360
rect 49974 38528 50030 38584
rect 50004 38106 50060 38108
rect 50084 38106 50140 38108
rect 50164 38106 50220 38108
rect 50244 38106 50300 38108
rect 50004 38054 50050 38106
rect 50050 38054 50060 38106
rect 50084 38054 50114 38106
rect 50114 38054 50126 38106
rect 50126 38054 50140 38106
rect 50164 38054 50178 38106
rect 50178 38054 50190 38106
rect 50190 38054 50220 38106
rect 50244 38054 50254 38106
rect 50254 38054 50300 38106
rect 50004 38052 50060 38054
rect 50084 38052 50140 38054
rect 50164 38052 50220 38054
rect 50244 38052 50300 38054
rect 50924 38650 50980 38652
rect 51004 38650 51060 38652
rect 51084 38650 51140 38652
rect 51164 38650 51220 38652
rect 50924 38598 50970 38650
rect 50970 38598 50980 38650
rect 51004 38598 51034 38650
rect 51034 38598 51046 38650
rect 51046 38598 51060 38650
rect 51084 38598 51098 38650
rect 51098 38598 51110 38650
rect 51110 38598 51140 38650
rect 51164 38598 51174 38650
rect 51174 38598 51220 38650
rect 50924 38596 50980 38598
rect 51004 38596 51060 38598
rect 51084 38596 51140 38598
rect 51164 38596 51220 38598
rect 50924 37562 50980 37564
rect 51004 37562 51060 37564
rect 51084 37562 51140 37564
rect 51164 37562 51220 37564
rect 50924 37510 50970 37562
rect 50970 37510 50980 37562
rect 51004 37510 51034 37562
rect 51034 37510 51046 37562
rect 51046 37510 51060 37562
rect 51084 37510 51098 37562
rect 51098 37510 51110 37562
rect 51110 37510 51140 37562
rect 51164 37510 51174 37562
rect 51174 37510 51220 37562
rect 50924 37508 50980 37510
rect 51004 37508 51060 37510
rect 51084 37508 51140 37510
rect 51164 37508 51220 37510
rect 52550 39480 52606 39536
rect 52826 39516 52828 39536
rect 52828 39516 52880 39536
rect 52880 39516 52882 39536
rect 52826 39480 52882 39516
rect 52090 38800 52146 38856
rect 58070 42200 58126 42256
rect 50004 37018 50060 37020
rect 50084 37018 50140 37020
rect 50164 37018 50220 37020
rect 50244 37018 50300 37020
rect 50004 36966 50050 37018
rect 50050 36966 50060 37018
rect 50084 36966 50114 37018
rect 50114 36966 50126 37018
rect 50126 36966 50140 37018
rect 50164 36966 50178 37018
rect 50178 36966 50190 37018
rect 50190 36966 50220 37018
rect 50244 36966 50254 37018
rect 50254 36966 50300 37018
rect 50004 36964 50060 36966
rect 50084 36964 50140 36966
rect 50164 36964 50220 36966
rect 50244 36964 50300 36966
rect 41694 36624 41750 36680
rect 55770 40976 55826 41032
rect 55218 38412 55274 38448
rect 55218 38392 55220 38412
rect 55220 38392 55272 38412
rect 55272 38392 55274 38412
rect 53838 37304 53894 37360
rect 56598 40996 56654 41032
rect 56598 40976 56600 40996
rect 56600 40976 56652 40996
rect 56652 40976 56654 40996
rect 42706 36352 42762 36408
rect 40130 35808 40186 35864
rect 30010 35672 30066 35728
rect 31022 35672 31078 35728
rect 33138 35672 33194 35728
rect 43534 35808 43590 35864
rect 56690 37848 56746 37904
rect 60738 41520 60794 41576
rect 62670 40024 62726 40080
rect 33598 35708 33600 35728
rect 33600 35708 33652 35728
rect 33652 35708 33654 35728
rect 33598 35672 33654 35708
rect 40038 35672 40094 35728
rect 42706 35672 42762 35728
rect 56046 35672 56102 35728
rect 62578 34992 62634 35048
rect 62762 36216 62818 36272
rect 62670 30882 62726 30938
rect 62762 29182 62818 29238
rect 62578 17176 62634 17232
rect 48962 1808 49018 1864
rect 49606 1808 49662 1864
rect 49698 1672 49754 1728
rect 63590 41112 63646 41168
rect 63314 36488 63370 36544
rect 63498 36080 63554 36136
rect 64694 39344 64750 39400
rect 63590 35536 63646 35592
rect 63498 33088 63554 33144
rect 63774 35944 63830 36000
rect 63866 35672 63922 35728
rect 62762 1400 62818 1456
rect 64344 37018 64400 37020
rect 64424 37018 64480 37020
rect 64504 37018 64560 37020
rect 64584 37018 64640 37020
rect 64344 36966 64390 37018
rect 64390 36966 64400 37018
rect 64424 36966 64454 37018
rect 64454 36966 64466 37018
rect 64466 36966 64480 37018
rect 64504 36966 64518 37018
rect 64518 36966 64530 37018
rect 64530 36966 64560 37018
rect 64584 36966 64594 37018
rect 64594 36966 64640 37018
rect 64344 36964 64400 36966
rect 64424 36964 64480 36966
rect 64504 36964 64560 36966
rect 64584 36964 64640 36966
rect 64344 35930 64400 35932
rect 64424 35930 64480 35932
rect 64504 35930 64560 35932
rect 64584 35930 64640 35932
rect 64344 35878 64390 35930
rect 64390 35878 64400 35930
rect 64424 35878 64454 35930
rect 64454 35878 64466 35930
rect 64466 35878 64480 35930
rect 64504 35878 64518 35930
rect 64518 35878 64530 35930
rect 64530 35878 64560 35930
rect 64584 35878 64594 35930
rect 64594 35878 64640 35930
rect 64344 35876 64400 35878
rect 64424 35876 64480 35878
rect 64504 35876 64560 35878
rect 64584 35876 64640 35878
rect 64344 34842 64400 34844
rect 64424 34842 64480 34844
rect 64504 34842 64560 34844
rect 64584 34842 64640 34844
rect 64344 34790 64390 34842
rect 64390 34790 64400 34842
rect 64424 34790 64454 34842
rect 64454 34790 64466 34842
rect 64466 34790 64480 34842
rect 64504 34790 64518 34842
rect 64518 34790 64530 34842
rect 64530 34790 64560 34842
rect 64584 34790 64594 34842
rect 64594 34790 64640 34842
rect 64344 34788 64400 34790
rect 64424 34788 64480 34790
rect 64504 34788 64560 34790
rect 64584 34788 64640 34790
rect 64344 33754 64400 33756
rect 64424 33754 64480 33756
rect 64504 33754 64560 33756
rect 64584 33754 64640 33756
rect 64344 33702 64390 33754
rect 64390 33702 64400 33754
rect 64424 33702 64454 33754
rect 64454 33702 64466 33754
rect 64466 33702 64480 33754
rect 64504 33702 64518 33754
rect 64518 33702 64530 33754
rect 64530 33702 64560 33754
rect 64584 33702 64594 33754
rect 64594 33702 64640 33754
rect 64344 33700 64400 33702
rect 64424 33700 64480 33702
rect 64504 33700 64560 33702
rect 64584 33700 64640 33702
rect 64344 32666 64400 32668
rect 64424 32666 64480 32668
rect 64504 32666 64560 32668
rect 64584 32666 64640 32668
rect 64344 32614 64390 32666
rect 64390 32614 64400 32666
rect 64424 32614 64454 32666
rect 64454 32614 64466 32666
rect 64466 32614 64480 32666
rect 64504 32614 64518 32666
rect 64518 32614 64530 32666
rect 64530 32614 64560 32666
rect 64584 32614 64594 32666
rect 64594 32614 64640 32666
rect 64344 32612 64400 32614
rect 64424 32612 64480 32614
rect 64504 32612 64560 32614
rect 64584 32612 64640 32614
rect 64694 32408 64750 32464
rect 64344 31578 64400 31580
rect 64424 31578 64480 31580
rect 64504 31578 64560 31580
rect 64584 31578 64640 31580
rect 64344 31526 64390 31578
rect 64390 31526 64400 31578
rect 64424 31526 64454 31578
rect 64454 31526 64466 31578
rect 64466 31526 64480 31578
rect 64504 31526 64518 31578
rect 64518 31526 64530 31578
rect 64530 31526 64560 31578
rect 64584 31526 64594 31578
rect 64594 31526 64640 31578
rect 64344 31524 64400 31526
rect 64424 31524 64480 31526
rect 64504 31524 64560 31526
rect 64584 31524 64640 31526
rect 64344 30490 64400 30492
rect 64424 30490 64480 30492
rect 64504 30490 64560 30492
rect 64584 30490 64640 30492
rect 64344 30438 64390 30490
rect 64390 30438 64400 30490
rect 64424 30438 64454 30490
rect 64454 30438 64466 30490
rect 64466 30438 64480 30490
rect 64504 30438 64518 30490
rect 64518 30438 64530 30490
rect 64530 30438 64560 30490
rect 64584 30438 64594 30490
rect 64594 30438 64640 30490
rect 64344 30436 64400 30438
rect 64424 30436 64480 30438
rect 64504 30436 64560 30438
rect 64584 30436 64640 30438
rect 64344 29402 64400 29404
rect 64424 29402 64480 29404
rect 64504 29402 64560 29404
rect 64584 29402 64640 29404
rect 64344 29350 64390 29402
rect 64390 29350 64400 29402
rect 64424 29350 64454 29402
rect 64454 29350 64466 29402
rect 64466 29350 64480 29402
rect 64504 29350 64518 29402
rect 64518 29350 64530 29402
rect 64530 29350 64560 29402
rect 64584 29350 64594 29402
rect 64594 29350 64640 29402
rect 64344 29348 64400 29350
rect 64424 29348 64480 29350
rect 64504 29348 64560 29350
rect 64584 29348 64640 29350
rect 64344 28314 64400 28316
rect 64424 28314 64480 28316
rect 64504 28314 64560 28316
rect 64584 28314 64640 28316
rect 64344 28262 64390 28314
rect 64390 28262 64400 28314
rect 64424 28262 64454 28314
rect 64454 28262 64466 28314
rect 64466 28262 64480 28314
rect 64504 28262 64518 28314
rect 64518 28262 64530 28314
rect 64530 28262 64560 28314
rect 64584 28262 64594 28314
rect 64594 28262 64640 28314
rect 64344 28260 64400 28262
rect 64424 28260 64480 28262
rect 64504 28260 64560 28262
rect 64584 28260 64640 28262
rect 64344 27226 64400 27228
rect 64424 27226 64480 27228
rect 64504 27226 64560 27228
rect 64584 27226 64640 27228
rect 64344 27174 64390 27226
rect 64390 27174 64400 27226
rect 64424 27174 64454 27226
rect 64454 27174 64466 27226
rect 64466 27174 64480 27226
rect 64504 27174 64518 27226
rect 64518 27174 64530 27226
rect 64530 27174 64560 27226
rect 64584 27174 64594 27226
rect 64594 27174 64640 27226
rect 64344 27172 64400 27174
rect 64424 27172 64480 27174
rect 64504 27172 64560 27174
rect 64584 27172 64640 27174
rect 64344 26138 64400 26140
rect 64424 26138 64480 26140
rect 64504 26138 64560 26140
rect 64584 26138 64640 26140
rect 64344 26086 64390 26138
rect 64390 26086 64400 26138
rect 64424 26086 64454 26138
rect 64454 26086 64466 26138
rect 64466 26086 64480 26138
rect 64504 26086 64518 26138
rect 64518 26086 64530 26138
rect 64530 26086 64560 26138
rect 64584 26086 64594 26138
rect 64594 26086 64640 26138
rect 64344 26084 64400 26086
rect 64424 26084 64480 26086
rect 64504 26084 64560 26086
rect 64584 26084 64640 26086
rect 64344 25050 64400 25052
rect 64424 25050 64480 25052
rect 64504 25050 64560 25052
rect 64584 25050 64640 25052
rect 64344 24998 64390 25050
rect 64390 24998 64400 25050
rect 64424 24998 64454 25050
rect 64454 24998 64466 25050
rect 64466 24998 64480 25050
rect 64504 24998 64518 25050
rect 64518 24998 64530 25050
rect 64530 24998 64560 25050
rect 64584 24998 64594 25050
rect 64594 24998 64640 25050
rect 64344 24996 64400 24998
rect 64424 24996 64480 24998
rect 64504 24996 64560 24998
rect 64584 24996 64640 24998
rect 64344 23962 64400 23964
rect 64424 23962 64480 23964
rect 64504 23962 64560 23964
rect 64584 23962 64640 23964
rect 64344 23910 64390 23962
rect 64390 23910 64400 23962
rect 64424 23910 64454 23962
rect 64454 23910 64466 23962
rect 64466 23910 64480 23962
rect 64504 23910 64518 23962
rect 64518 23910 64530 23962
rect 64530 23910 64560 23962
rect 64584 23910 64594 23962
rect 64594 23910 64640 23962
rect 64344 23908 64400 23910
rect 64424 23908 64480 23910
rect 64504 23908 64560 23910
rect 64584 23908 64640 23910
rect 64344 22874 64400 22876
rect 64424 22874 64480 22876
rect 64504 22874 64560 22876
rect 64584 22874 64640 22876
rect 64344 22822 64390 22874
rect 64390 22822 64400 22874
rect 64424 22822 64454 22874
rect 64454 22822 64466 22874
rect 64466 22822 64480 22874
rect 64504 22822 64518 22874
rect 64518 22822 64530 22874
rect 64530 22822 64560 22874
rect 64584 22822 64594 22874
rect 64594 22822 64640 22874
rect 64344 22820 64400 22822
rect 64424 22820 64480 22822
rect 64504 22820 64560 22822
rect 64584 22820 64640 22822
rect 64970 31748 65026 31784
rect 64970 31728 64972 31748
rect 64972 31728 65024 31748
rect 65024 31728 65026 31748
rect 65264 37562 65320 37564
rect 65344 37562 65400 37564
rect 65424 37562 65480 37564
rect 65504 37562 65560 37564
rect 65264 37510 65310 37562
rect 65310 37510 65320 37562
rect 65344 37510 65374 37562
rect 65374 37510 65386 37562
rect 65386 37510 65400 37562
rect 65424 37510 65438 37562
rect 65438 37510 65450 37562
rect 65450 37510 65480 37562
rect 65504 37510 65514 37562
rect 65514 37510 65560 37562
rect 65264 37508 65320 37510
rect 65344 37508 65400 37510
rect 65424 37508 65480 37510
rect 65504 37508 65560 37510
rect 65614 36624 65670 36680
rect 65264 36474 65320 36476
rect 65344 36474 65400 36476
rect 65424 36474 65480 36476
rect 65504 36474 65560 36476
rect 65264 36422 65310 36474
rect 65310 36422 65320 36474
rect 65344 36422 65374 36474
rect 65374 36422 65386 36474
rect 65386 36422 65400 36474
rect 65424 36422 65438 36474
rect 65438 36422 65450 36474
rect 65450 36422 65480 36474
rect 65504 36422 65514 36474
rect 65514 36422 65560 36474
rect 65264 36420 65320 36422
rect 65344 36420 65400 36422
rect 65424 36420 65480 36422
rect 65504 36420 65560 36422
rect 65264 35386 65320 35388
rect 65344 35386 65400 35388
rect 65424 35386 65480 35388
rect 65504 35386 65560 35388
rect 65264 35334 65310 35386
rect 65310 35334 65320 35386
rect 65344 35334 65374 35386
rect 65374 35334 65386 35386
rect 65386 35334 65400 35386
rect 65424 35334 65438 35386
rect 65438 35334 65450 35386
rect 65450 35334 65480 35386
rect 65504 35334 65514 35386
rect 65514 35334 65560 35386
rect 65264 35332 65320 35334
rect 65344 35332 65400 35334
rect 65424 35332 65480 35334
rect 65504 35332 65560 35334
rect 65264 34298 65320 34300
rect 65344 34298 65400 34300
rect 65424 34298 65480 34300
rect 65504 34298 65560 34300
rect 65264 34246 65310 34298
rect 65310 34246 65320 34298
rect 65344 34246 65374 34298
rect 65374 34246 65386 34298
rect 65386 34246 65400 34298
rect 65424 34246 65438 34298
rect 65438 34246 65450 34298
rect 65450 34246 65480 34298
rect 65504 34246 65514 34298
rect 65514 34246 65560 34298
rect 65264 34244 65320 34246
rect 65344 34244 65400 34246
rect 65424 34244 65480 34246
rect 65504 34244 65560 34246
rect 65264 33210 65320 33212
rect 65344 33210 65400 33212
rect 65424 33210 65480 33212
rect 65504 33210 65560 33212
rect 65264 33158 65310 33210
rect 65310 33158 65320 33210
rect 65344 33158 65374 33210
rect 65374 33158 65386 33210
rect 65386 33158 65400 33210
rect 65424 33158 65438 33210
rect 65438 33158 65450 33210
rect 65450 33158 65480 33210
rect 65504 33158 65514 33210
rect 65514 33158 65560 33210
rect 65264 33156 65320 33158
rect 65344 33156 65400 33158
rect 65424 33156 65480 33158
rect 65504 33156 65560 33158
rect 65264 32122 65320 32124
rect 65344 32122 65400 32124
rect 65424 32122 65480 32124
rect 65504 32122 65560 32124
rect 65264 32070 65310 32122
rect 65310 32070 65320 32122
rect 65344 32070 65374 32122
rect 65374 32070 65386 32122
rect 65386 32070 65400 32122
rect 65424 32070 65438 32122
rect 65438 32070 65450 32122
rect 65450 32070 65480 32122
rect 65504 32070 65514 32122
rect 65514 32070 65560 32122
rect 65264 32068 65320 32070
rect 65344 32068 65400 32070
rect 65424 32068 65480 32070
rect 65504 32068 65560 32070
rect 65338 31728 65394 31784
rect 65264 31034 65320 31036
rect 65344 31034 65400 31036
rect 65424 31034 65480 31036
rect 65504 31034 65560 31036
rect 65264 30982 65310 31034
rect 65310 30982 65320 31034
rect 65344 30982 65374 31034
rect 65374 30982 65386 31034
rect 65386 30982 65400 31034
rect 65424 30982 65438 31034
rect 65438 30982 65450 31034
rect 65450 30982 65480 31034
rect 65504 30982 65514 31034
rect 65514 30982 65560 31034
rect 65264 30980 65320 30982
rect 65344 30980 65400 30982
rect 65424 30980 65480 30982
rect 65504 30980 65560 30982
rect 65264 29946 65320 29948
rect 65344 29946 65400 29948
rect 65424 29946 65480 29948
rect 65504 29946 65560 29948
rect 65264 29894 65310 29946
rect 65310 29894 65320 29946
rect 65344 29894 65374 29946
rect 65374 29894 65386 29946
rect 65386 29894 65400 29946
rect 65424 29894 65438 29946
rect 65438 29894 65450 29946
rect 65450 29894 65480 29946
rect 65504 29894 65514 29946
rect 65514 29894 65560 29946
rect 65264 29892 65320 29894
rect 65344 29892 65400 29894
rect 65424 29892 65480 29894
rect 65504 29892 65560 29894
rect 65890 31728 65946 31784
rect 65264 28858 65320 28860
rect 65344 28858 65400 28860
rect 65424 28858 65480 28860
rect 65504 28858 65560 28860
rect 65264 28806 65310 28858
rect 65310 28806 65320 28858
rect 65344 28806 65374 28858
rect 65374 28806 65386 28858
rect 65386 28806 65400 28858
rect 65424 28806 65438 28858
rect 65438 28806 65450 28858
rect 65450 28806 65480 28858
rect 65504 28806 65514 28858
rect 65514 28806 65560 28858
rect 65264 28804 65320 28806
rect 65344 28804 65400 28806
rect 65424 28804 65480 28806
rect 65504 28804 65560 28806
rect 65264 27770 65320 27772
rect 65344 27770 65400 27772
rect 65424 27770 65480 27772
rect 65504 27770 65560 27772
rect 65264 27718 65310 27770
rect 65310 27718 65320 27770
rect 65344 27718 65374 27770
rect 65374 27718 65386 27770
rect 65386 27718 65400 27770
rect 65424 27718 65438 27770
rect 65438 27718 65450 27770
rect 65450 27718 65480 27770
rect 65504 27718 65514 27770
rect 65514 27718 65560 27770
rect 65264 27716 65320 27718
rect 65344 27716 65400 27718
rect 65424 27716 65480 27718
rect 65504 27716 65560 27718
rect 65264 26682 65320 26684
rect 65344 26682 65400 26684
rect 65424 26682 65480 26684
rect 65504 26682 65560 26684
rect 65264 26630 65310 26682
rect 65310 26630 65320 26682
rect 65344 26630 65374 26682
rect 65374 26630 65386 26682
rect 65386 26630 65400 26682
rect 65424 26630 65438 26682
rect 65438 26630 65450 26682
rect 65450 26630 65480 26682
rect 65504 26630 65514 26682
rect 65514 26630 65560 26682
rect 65264 26628 65320 26630
rect 65344 26628 65400 26630
rect 65424 26628 65480 26630
rect 65504 26628 65560 26630
rect 65264 25594 65320 25596
rect 65344 25594 65400 25596
rect 65424 25594 65480 25596
rect 65504 25594 65560 25596
rect 65264 25542 65310 25594
rect 65310 25542 65320 25594
rect 65344 25542 65374 25594
rect 65374 25542 65386 25594
rect 65386 25542 65400 25594
rect 65424 25542 65438 25594
rect 65438 25542 65450 25594
rect 65450 25542 65480 25594
rect 65504 25542 65514 25594
rect 65514 25542 65560 25594
rect 65264 25540 65320 25542
rect 65344 25540 65400 25542
rect 65424 25540 65480 25542
rect 65504 25540 65560 25542
rect 65264 24506 65320 24508
rect 65344 24506 65400 24508
rect 65424 24506 65480 24508
rect 65504 24506 65560 24508
rect 65264 24454 65310 24506
rect 65310 24454 65320 24506
rect 65344 24454 65374 24506
rect 65374 24454 65386 24506
rect 65386 24454 65400 24506
rect 65424 24454 65438 24506
rect 65438 24454 65450 24506
rect 65450 24454 65480 24506
rect 65504 24454 65514 24506
rect 65514 24454 65560 24506
rect 65264 24452 65320 24454
rect 65344 24452 65400 24454
rect 65424 24452 65480 24454
rect 65504 24452 65560 24454
rect 65264 23418 65320 23420
rect 65344 23418 65400 23420
rect 65424 23418 65480 23420
rect 65504 23418 65560 23420
rect 65264 23366 65310 23418
rect 65310 23366 65320 23418
rect 65344 23366 65374 23418
rect 65374 23366 65386 23418
rect 65386 23366 65400 23418
rect 65424 23366 65438 23418
rect 65438 23366 65450 23418
rect 65450 23366 65480 23418
rect 65504 23366 65514 23418
rect 65514 23366 65560 23418
rect 65264 23364 65320 23366
rect 65344 23364 65400 23366
rect 65424 23364 65480 23366
rect 65504 23364 65560 23366
rect 64344 21786 64400 21788
rect 64424 21786 64480 21788
rect 64504 21786 64560 21788
rect 64584 21786 64640 21788
rect 64344 21734 64390 21786
rect 64390 21734 64400 21786
rect 64424 21734 64454 21786
rect 64454 21734 64466 21786
rect 64466 21734 64480 21786
rect 64504 21734 64518 21786
rect 64518 21734 64530 21786
rect 64530 21734 64560 21786
rect 64584 21734 64594 21786
rect 64594 21734 64640 21786
rect 64344 21732 64400 21734
rect 64424 21732 64480 21734
rect 64504 21732 64560 21734
rect 64584 21732 64640 21734
rect 64344 20698 64400 20700
rect 64424 20698 64480 20700
rect 64504 20698 64560 20700
rect 64584 20698 64640 20700
rect 64344 20646 64390 20698
rect 64390 20646 64400 20698
rect 64424 20646 64454 20698
rect 64454 20646 64466 20698
rect 64466 20646 64480 20698
rect 64504 20646 64518 20698
rect 64518 20646 64530 20698
rect 64530 20646 64560 20698
rect 64584 20646 64594 20698
rect 64594 20646 64640 20698
rect 64344 20644 64400 20646
rect 64424 20644 64480 20646
rect 64504 20644 64560 20646
rect 64584 20644 64640 20646
rect 65264 22330 65320 22332
rect 65344 22330 65400 22332
rect 65424 22330 65480 22332
rect 65504 22330 65560 22332
rect 65264 22278 65310 22330
rect 65310 22278 65320 22330
rect 65344 22278 65374 22330
rect 65374 22278 65386 22330
rect 65386 22278 65400 22330
rect 65424 22278 65438 22330
rect 65438 22278 65450 22330
rect 65450 22278 65480 22330
rect 65504 22278 65514 22330
rect 65514 22278 65560 22330
rect 65264 22276 65320 22278
rect 65344 22276 65400 22278
rect 65424 22276 65480 22278
rect 65504 22276 65560 22278
rect 65264 21242 65320 21244
rect 65344 21242 65400 21244
rect 65424 21242 65480 21244
rect 65504 21242 65560 21244
rect 65264 21190 65310 21242
rect 65310 21190 65320 21242
rect 65344 21190 65374 21242
rect 65374 21190 65386 21242
rect 65386 21190 65400 21242
rect 65424 21190 65438 21242
rect 65438 21190 65450 21242
rect 65450 21190 65480 21242
rect 65504 21190 65514 21242
rect 65514 21190 65560 21242
rect 65264 21188 65320 21190
rect 65344 21188 65400 21190
rect 65424 21188 65480 21190
rect 65504 21188 65560 21190
rect 64344 19610 64400 19612
rect 64424 19610 64480 19612
rect 64504 19610 64560 19612
rect 64584 19610 64640 19612
rect 64344 19558 64390 19610
rect 64390 19558 64400 19610
rect 64424 19558 64454 19610
rect 64454 19558 64466 19610
rect 64466 19558 64480 19610
rect 64504 19558 64518 19610
rect 64518 19558 64530 19610
rect 64530 19558 64560 19610
rect 64584 19558 64594 19610
rect 64594 19558 64640 19610
rect 64344 19556 64400 19558
rect 64424 19556 64480 19558
rect 64504 19556 64560 19558
rect 64584 19556 64640 19558
rect 64344 18522 64400 18524
rect 64424 18522 64480 18524
rect 64504 18522 64560 18524
rect 64584 18522 64640 18524
rect 64344 18470 64390 18522
rect 64390 18470 64400 18522
rect 64424 18470 64454 18522
rect 64454 18470 64466 18522
rect 64466 18470 64480 18522
rect 64504 18470 64518 18522
rect 64518 18470 64530 18522
rect 64530 18470 64560 18522
rect 64584 18470 64594 18522
rect 64594 18470 64640 18522
rect 64344 18468 64400 18470
rect 64424 18468 64480 18470
rect 64504 18468 64560 18470
rect 64584 18468 64640 18470
rect 64694 17856 64750 17912
rect 64344 17434 64400 17436
rect 64424 17434 64480 17436
rect 64504 17434 64560 17436
rect 64584 17434 64640 17436
rect 64344 17382 64390 17434
rect 64390 17382 64400 17434
rect 64424 17382 64454 17434
rect 64454 17382 64466 17434
rect 64466 17382 64480 17434
rect 64504 17382 64518 17434
rect 64518 17382 64530 17434
rect 64530 17382 64560 17434
rect 64584 17382 64594 17434
rect 64594 17382 64640 17434
rect 64344 17380 64400 17382
rect 64424 17380 64480 17382
rect 64504 17380 64560 17382
rect 64584 17380 64640 17382
rect 64344 16346 64400 16348
rect 64424 16346 64480 16348
rect 64504 16346 64560 16348
rect 64584 16346 64640 16348
rect 64344 16294 64390 16346
rect 64390 16294 64400 16346
rect 64424 16294 64454 16346
rect 64454 16294 64466 16346
rect 64466 16294 64480 16346
rect 64504 16294 64518 16346
rect 64518 16294 64530 16346
rect 64530 16294 64560 16346
rect 64584 16294 64594 16346
rect 64594 16294 64640 16346
rect 64344 16292 64400 16294
rect 64424 16292 64480 16294
rect 64504 16292 64560 16294
rect 64584 16292 64640 16294
rect 65264 20154 65320 20156
rect 65344 20154 65400 20156
rect 65424 20154 65480 20156
rect 65504 20154 65560 20156
rect 65264 20102 65310 20154
rect 65310 20102 65320 20154
rect 65344 20102 65374 20154
rect 65374 20102 65386 20154
rect 65386 20102 65400 20154
rect 65424 20102 65438 20154
rect 65438 20102 65450 20154
rect 65450 20102 65480 20154
rect 65504 20102 65514 20154
rect 65514 20102 65560 20154
rect 65264 20100 65320 20102
rect 65344 20100 65400 20102
rect 65424 20100 65480 20102
rect 65504 20100 65560 20102
rect 65264 19066 65320 19068
rect 65344 19066 65400 19068
rect 65424 19066 65480 19068
rect 65504 19066 65560 19068
rect 65264 19014 65310 19066
rect 65310 19014 65320 19066
rect 65344 19014 65374 19066
rect 65374 19014 65386 19066
rect 65386 19014 65400 19066
rect 65424 19014 65438 19066
rect 65438 19014 65450 19066
rect 65450 19014 65480 19066
rect 65504 19014 65514 19066
rect 65514 19014 65560 19066
rect 65264 19012 65320 19014
rect 65344 19012 65400 19014
rect 65424 19012 65480 19014
rect 65504 19012 65560 19014
rect 64344 15258 64400 15260
rect 64424 15258 64480 15260
rect 64504 15258 64560 15260
rect 64584 15258 64640 15260
rect 64344 15206 64390 15258
rect 64390 15206 64400 15258
rect 64424 15206 64454 15258
rect 64454 15206 64466 15258
rect 64466 15206 64480 15258
rect 64504 15206 64518 15258
rect 64518 15206 64530 15258
rect 64530 15206 64560 15258
rect 64584 15206 64594 15258
rect 64594 15206 64640 15258
rect 64344 15204 64400 15206
rect 64424 15204 64480 15206
rect 64504 15204 64560 15206
rect 64584 15204 64640 15206
rect 64344 14170 64400 14172
rect 64424 14170 64480 14172
rect 64504 14170 64560 14172
rect 64584 14170 64640 14172
rect 64344 14118 64390 14170
rect 64390 14118 64400 14170
rect 64424 14118 64454 14170
rect 64454 14118 64466 14170
rect 64466 14118 64480 14170
rect 64504 14118 64518 14170
rect 64518 14118 64530 14170
rect 64530 14118 64560 14170
rect 64584 14118 64594 14170
rect 64594 14118 64640 14170
rect 64344 14116 64400 14118
rect 64424 14116 64480 14118
rect 64504 14116 64560 14118
rect 64584 14116 64640 14118
rect 64344 13082 64400 13084
rect 64424 13082 64480 13084
rect 64504 13082 64560 13084
rect 64584 13082 64640 13084
rect 64344 13030 64390 13082
rect 64390 13030 64400 13082
rect 64424 13030 64454 13082
rect 64454 13030 64466 13082
rect 64466 13030 64480 13082
rect 64504 13030 64518 13082
rect 64518 13030 64530 13082
rect 64530 13030 64560 13082
rect 64584 13030 64594 13082
rect 64594 13030 64640 13082
rect 64344 13028 64400 13030
rect 64424 13028 64480 13030
rect 64504 13028 64560 13030
rect 64584 13028 64640 13030
rect 64786 15700 64842 15736
rect 64786 15680 64788 15700
rect 64788 15680 64840 15700
rect 64840 15680 64842 15700
rect 65264 17978 65320 17980
rect 65344 17978 65400 17980
rect 65424 17978 65480 17980
rect 65504 17978 65560 17980
rect 65264 17926 65310 17978
rect 65310 17926 65320 17978
rect 65344 17926 65374 17978
rect 65374 17926 65386 17978
rect 65386 17926 65400 17978
rect 65424 17926 65438 17978
rect 65438 17926 65450 17978
rect 65450 17926 65480 17978
rect 65504 17926 65514 17978
rect 65514 17926 65560 17978
rect 65264 17924 65320 17926
rect 65344 17924 65400 17926
rect 65424 17924 65480 17926
rect 65504 17924 65560 17926
rect 65264 16890 65320 16892
rect 65344 16890 65400 16892
rect 65424 16890 65480 16892
rect 65504 16890 65560 16892
rect 65264 16838 65310 16890
rect 65310 16838 65320 16890
rect 65344 16838 65374 16890
rect 65374 16838 65386 16890
rect 65386 16838 65400 16890
rect 65424 16838 65438 16890
rect 65438 16838 65450 16890
rect 65450 16838 65480 16890
rect 65504 16838 65514 16890
rect 65514 16838 65560 16890
rect 65264 16836 65320 16838
rect 65344 16836 65400 16838
rect 65424 16836 65480 16838
rect 65504 16836 65560 16838
rect 65264 15802 65320 15804
rect 65344 15802 65400 15804
rect 65424 15802 65480 15804
rect 65504 15802 65560 15804
rect 65264 15750 65310 15802
rect 65310 15750 65320 15802
rect 65344 15750 65374 15802
rect 65374 15750 65386 15802
rect 65386 15750 65400 15802
rect 65424 15750 65438 15802
rect 65438 15750 65450 15802
rect 65450 15750 65480 15802
rect 65504 15750 65514 15802
rect 65514 15750 65560 15802
rect 65264 15748 65320 15750
rect 65344 15748 65400 15750
rect 65424 15748 65480 15750
rect 65504 15748 65560 15750
rect 64344 11994 64400 11996
rect 64424 11994 64480 11996
rect 64504 11994 64560 11996
rect 64584 11994 64640 11996
rect 64344 11942 64390 11994
rect 64390 11942 64400 11994
rect 64424 11942 64454 11994
rect 64454 11942 64466 11994
rect 64466 11942 64480 11994
rect 64504 11942 64518 11994
rect 64518 11942 64530 11994
rect 64530 11942 64560 11994
rect 64584 11942 64594 11994
rect 64594 11942 64640 11994
rect 64344 11940 64400 11942
rect 64424 11940 64480 11942
rect 64504 11940 64560 11942
rect 64584 11940 64640 11942
rect 64344 10906 64400 10908
rect 64424 10906 64480 10908
rect 64504 10906 64560 10908
rect 64584 10906 64640 10908
rect 64344 10854 64390 10906
rect 64390 10854 64400 10906
rect 64424 10854 64454 10906
rect 64454 10854 64466 10906
rect 64466 10854 64480 10906
rect 64504 10854 64518 10906
rect 64518 10854 64530 10906
rect 64530 10854 64560 10906
rect 64584 10854 64594 10906
rect 64594 10854 64640 10906
rect 64344 10852 64400 10854
rect 64424 10852 64480 10854
rect 64504 10852 64560 10854
rect 64584 10852 64640 10854
rect 65264 14714 65320 14716
rect 65344 14714 65400 14716
rect 65424 14714 65480 14716
rect 65504 14714 65560 14716
rect 65264 14662 65310 14714
rect 65310 14662 65320 14714
rect 65344 14662 65374 14714
rect 65374 14662 65386 14714
rect 65386 14662 65400 14714
rect 65424 14662 65438 14714
rect 65438 14662 65450 14714
rect 65450 14662 65480 14714
rect 65504 14662 65514 14714
rect 65514 14662 65560 14714
rect 65264 14660 65320 14662
rect 65344 14660 65400 14662
rect 65424 14660 65480 14662
rect 65504 14660 65560 14662
rect 65264 13626 65320 13628
rect 65344 13626 65400 13628
rect 65424 13626 65480 13628
rect 65504 13626 65560 13628
rect 65264 13574 65310 13626
rect 65310 13574 65320 13626
rect 65344 13574 65374 13626
rect 65374 13574 65386 13626
rect 65386 13574 65400 13626
rect 65424 13574 65438 13626
rect 65438 13574 65450 13626
rect 65450 13574 65480 13626
rect 65504 13574 65514 13626
rect 65514 13574 65560 13626
rect 65264 13572 65320 13574
rect 65344 13572 65400 13574
rect 65424 13572 65480 13574
rect 65504 13572 65560 13574
rect 65264 12538 65320 12540
rect 65344 12538 65400 12540
rect 65424 12538 65480 12540
rect 65504 12538 65560 12540
rect 65264 12486 65310 12538
rect 65310 12486 65320 12538
rect 65344 12486 65374 12538
rect 65374 12486 65386 12538
rect 65386 12486 65400 12538
rect 65424 12486 65438 12538
rect 65438 12486 65450 12538
rect 65450 12486 65480 12538
rect 65504 12486 65514 12538
rect 65514 12486 65560 12538
rect 65264 12484 65320 12486
rect 65344 12484 65400 12486
rect 65424 12484 65480 12486
rect 65504 12484 65560 12486
rect 65264 11450 65320 11452
rect 65344 11450 65400 11452
rect 65424 11450 65480 11452
rect 65504 11450 65560 11452
rect 65264 11398 65310 11450
rect 65310 11398 65320 11450
rect 65344 11398 65374 11450
rect 65374 11398 65386 11450
rect 65386 11398 65400 11450
rect 65424 11398 65438 11450
rect 65438 11398 65450 11450
rect 65450 11398 65480 11450
rect 65504 11398 65514 11450
rect 65514 11398 65560 11450
rect 65264 11396 65320 11398
rect 65344 11396 65400 11398
rect 65424 11396 65480 11398
rect 65504 11396 65560 11398
rect 64344 9818 64400 9820
rect 64424 9818 64480 9820
rect 64504 9818 64560 9820
rect 64584 9818 64640 9820
rect 64344 9766 64390 9818
rect 64390 9766 64400 9818
rect 64424 9766 64454 9818
rect 64454 9766 64466 9818
rect 64466 9766 64480 9818
rect 64504 9766 64518 9818
rect 64518 9766 64530 9818
rect 64530 9766 64560 9818
rect 64584 9766 64594 9818
rect 64594 9766 64640 9818
rect 64344 9764 64400 9766
rect 64424 9764 64480 9766
rect 64504 9764 64560 9766
rect 64584 9764 64640 9766
rect 65264 10362 65320 10364
rect 65344 10362 65400 10364
rect 65424 10362 65480 10364
rect 65504 10362 65560 10364
rect 65264 10310 65310 10362
rect 65310 10310 65320 10362
rect 65344 10310 65374 10362
rect 65374 10310 65386 10362
rect 65386 10310 65400 10362
rect 65424 10310 65438 10362
rect 65438 10310 65450 10362
rect 65450 10310 65480 10362
rect 65504 10310 65514 10362
rect 65514 10310 65560 10362
rect 65264 10308 65320 10310
rect 65344 10308 65400 10310
rect 65424 10308 65480 10310
rect 65504 10308 65560 10310
rect 64142 6840 64198 6896
rect 64344 8730 64400 8732
rect 64424 8730 64480 8732
rect 64504 8730 64560 8732
rect 64584 8730 64640 8732
rect 64344 8678 64390 8730
rect 64390 8678 64400 8730
rect 64424 8678 64454 8730
rect 64454 8678 64466 8730
rect 64466 8678 64480 8730
rect 64504 8678 64518 8730
rect 64518 8678 64530 8730
rect 64530 8678 64560 8730
rect 64584 8678 64594 8730
rect 64594 8678 64640 8730
rect 64344 8676 64400 8678
rect 64424 8676 64480 8678
rect 64504 8676 64560 8678
rect 64584 8676 64640 8678
rect 64344 7642 64400 7644
rect 64424 7642 64480 7644
rect 64504 7642 64560 7644
rect 64584 7642 64640 7644
rect 64344 7590 64390 7642
rect 64390 7590 64400 7642
rect 64424 7590 64454 7642
rect 64454 7590 64466 7642
rect 64466 7590 64480 7642
rect 64504 7590 64518 7642
rect 64518 7590 64530 7642
rect 64530 7590 64560 7642
rect 64584 7590 64594 7642
rect 64594 7590 64640 7642
rect 64344 7588 64400 7590
rect 64424 7588 64480 7590
rect 64504 7588 64560 7590
rect 64584 7588 64640 7590
rect 64510 7384 64566 7440
rect 64602 6860 64658 6896
rect 64602 6840 64604 6860
rect 64604 6840 64656 6860
rect 64656 6840 64658 6860
rect 64344 6554 64400 6556
rect 64424 6554 64480 6556
rect 64504 6554 64560 6556
rect 64584 6554 64640 6556
rect 64344 6502 64390 6554
rect 64390 6502 64400 6554
rect 64424 6502 64454 6554
rect 64454 6502 64466 6554
rect 64466 6502 64480 6554
rect 64504 6502 64518 6554
rect 64518 6502 64530 6554
rect 64530 6502 64560 6554
rect 64584 6502 64594 6554
rect 64594 6502 64640 6554
rect 64344 6500 64400 6502
rect 64424 6500 64480 6502
rect 64504 6500 64560 6502
rect 64584 6500 64640 6502
rect 64344 5466 64400 5468
rect 64424 5466 64480 5468
rect 64504 5466 64560 5468
rect 64584 5466 64640 5468
rect 64344 5414 64390 5466
rect 64390 5414 64400 5466
rect 64424 5414 64454 5466
rect 64454 5414 64466 5466
rect 64466 5414 64480 5466
rect 64504 5414 64518 5466
rect 64518 5414 64530 5466
rect 64530 5414 64560 5466
rect 64584 5414 64594 5466
rect 64594 5414 64640 5466
rect 64344 5412 64400 5414
rect 64424 5412 64480 5414
rect 64504 5412 64560 5414
rect 64584 5412 64640 5414
rect 65264 9274 65320 9276
rect 65344 9274 65400 9276
rect 65424 9274 65480 9276
rect 65504 9274 65560 9276
rect 65264 9222 65310 9274
rect 65310 9222 65320 9274
rect 65344 9222 65374 9274
rect 65374 9222 65386 9274
rect 65386 9222 65400 9274
rect 65424 9222 65438 9274
rect 65438 9222 65450 9274
rect 65450 9222 65480 9274
rect 65504 9222 65514 9274
rect 65514 9222 65560 9274
rect 65264 9220 65320 9222
rect 65344 9220 65400 9222
rect 65424 9220 65480 9222
rect 65504 9220 65560 9222
rect 66166 31864 66222 31920
rect 65264 8186 65320 8188
rect 65344 8186 65400 8188
rect 65424 8186 65480 8188
rect 65504 8186 65560 8188
rect 65264 8134 65310 8186
rect 65310 8134 65320 8186
rect 65344 8134 65374 8186
rect 65374 8134 65386 8186
rect 65386 8134 65400 8186
rect 65424 8134 65438 8186
rect 65438 8134 65450 8186
rect 65450 8134 65480 8186
rect 65504 8134 65514 8186
rect 65514 8134 65560 8186
rect 65264 8132 65320 8134
rect 65344 8132 65400 8134
rect 65424 8132 65480 8134
rect 65504 8132 65560 8134
rect 65264 7098 65320 7100
rect 65344 7098 65400 7100
rect 65424 7098 65480 7100
rect 65504 7098 65560 7100
rect 65264 7046 65310 7098
rect 65310 7046 65320 7098
rect 65344 7046 65374 7098
rect 65374 7046 65386 7098
rect 65386 7046 65400 7098
rect 65424 7046 65438 7098
rect 65438 7046 65450 7098
rect 65450 7046 65480 7098
rect 65504 7046 65514 7098
rect 65514 7046 65560 7098
rect 65264 7044 65320 7046
rect 65344 7044 65400 7046
rect 65424 7044 65480 7046
rect 65504 7044 65560 7046
rect 64344 4378 64400 4380
rect 64424 4378 64480 4380
rect 64504 4378 64560 4380
rect 64584 4378 64640 4380
rect 64344 4326 64390 4378
rect 64390 4326 64400 4378
rect 64424 4326 64454 4378
rect 64454 4326 64466 4378
rect 64466 4326 64480 4378
rect 64504 4326 64518 4378
rect 64518 4326 64530 4378
rect 64530 4326 64560 4378
rect 64584 4326 64594 4378
rect 64594 4326 64640 4378
rect 64344 4324 64400 4326
rect 64424 4324 64480 4326
rect 64504 4324 64560 4326
rect 64584 4324 64640 4326
rect 64344 3290 64400 3292
rect 64424 3290 64480 3292
rect 64504 3290 64560 3292
rect 64584 3290 64640 3292
rect 64344 3238 64390 3290
rect 64390 3238 64400 3290
rect 64424 3238 64454 3290
rect 64454 3238 64466 3290
rect 64466 3238 64480 3290
rect 64504 3238 64518 3290
rect 64518 3238 64530 3290
rect 64530 3238 64560 3290
rect 64584 3238 64594 3290
rect 64594 3238 64640 3290
rect 64344 3236 64400 3238
rect 64424 3236 64480 3238
rect 64504 3236 64560 3238
rect 64584 3236 64640 3238
rect 65264 6010 65320 6012
rect 65344 6010 65400 6012
rect 65424 6010 65480 6012
rect 65504 6010 65560 6012
rect 65264 5958 65310 6010
rect 65310 5958 65320 6010
rect 65344 5958 65374 6010
rect 65374 5958 65386 6010
rect 65386 5958 65400 6010
rect 65424 5958 65438 6010
rect 65438 5958 65450 6010
rect 65450 5958 65480 6010
rect 65504 5958 65514 6010
rect 65514 5958 65560 6010
rect 65264 5956 65320 5958
rect 65344 5956 65400 5958
rect 65424 5956 65480 5958
rect 65504 5956 65560 5958
rect 65264 4922 65320 4924
rect 65344 4922 65400 4924
rect 65424 4922 65480 4924
rect 65504 4922 65560 4924
rect 65264 4870 65310 4922
rect 65310 4870 65320 4922
rect 65344 4870 65374 4922
rect 65374 4870 65386 4922
rect 65386 4870 65400 4922
rect 65424 4870 65438 4922
rect 65438 4870 65450 4922
rect 65450 4870 65480 4922
rect 65504 4870 65514 4922
rect 65514 4870 65560 4922
rect 65264 4868 65320 4870
rect 65344 4868 65400 4870
rect 65424 4868 65480 4870
rect 65504 4868 65560 4870
rect 63682 1808 63738 1864
rect 64344 2202 64400 2204
rect 64424 2202 64480 2204
rect 64504 2202 64560 2204
rect 64584 2202 64640 2204
rect 64344 2150 64390 2202
rect 64390 2150 64400 2202
rect 64424 2150 64454 2202
rect 64454 2150 64466 2202
rect 64466 2150 64480 2202
rect 64504 2150 64518 2202
rect 64518 2150 64530 2202
rect 64530 2150 64560 2202
rect 64584 2150 64594 2202
rect 64594 2150 64640 2202
rect 64344 2148 64400 2150
rect 64424 2148 64480 2150
rect 64504 2148 64560 2150
rect 64584 2148 64640 2150
rect 65264 3834 65320 3836
rect 65344 3834 65400 3836
rect 65424 3834 65480 3836
rect 65504 3834 65560 3836
rect 65264 3782 65310 3834
rect 65310 3782 65320 3834
rect 65344 3782 65374 3834
rect 65374 3782 65386 3834
rect 65386 3782 65400 3834
rect 65424 3782 65438 3834
rect 65438 3782 65450 3834
rect 65450 3782 65480 3834
rect 65504 3782 65514 3834
rect 65514 3782 65560 3834
rect 65264 3780 65320 3782
rect 65344 3780 65400 3782
rect 65424 3780 65480 3782
rect 65504 3780 65560 3782
rect 65264 2746 65320 2748
rect 65344 2746 65400 2748
rect 65424 2746 65480 2748
rect 65504 2746 65560 2748
rect 65264 2694 65310 2746
rect 65310 2694 65320 2746
rect 65344 2694 65374 2746
rect 65374 2694 65386 2746
rect 65386 2694 65400 2746
rect 65424 2694 65438 2746
rect 65438 2694 65450 2746
rect 65450 2694 65480 2746
rect 65504 2694 65514 2746
rect 65514 2694 65560 2746
rect 65264 2692 65320 2694
rect 65344 2692 65400 2694
rect 65424 2692 65480 2694
rect 65504 2692 65560 2694
rect 65264 1658 65320 1660
rect 65344 1658 65400 1660
rect 65424 1658 65480 1660
rect 65504 1658 65560 1660
rect 65264 1606 65310 1658
rect 65310 1606 65320 1658
rect 65344 1606 65374 1658
rect 65374 1606 65386 1658
rect 65386 1606 65400 1658
rect 65424 1606 65438 1658
rect 65438 1606 65450 1658
rect 65450 1606 65480 1658
rect 65504 1606 65514 1658
rect 65514 1606 65560 1658
rect 65264 1604 65320 1606
rect 65344 1604 65400 1606
rect 65424 1604 65480 1606
rect 65504 1604 65560 1606
rect 62946 1264 63002 1320
rect 64344 1114 64400 1116
rect 64424 1114 64480 1116
rect 64504 1114 64560 1116
rect 64584 1114 64640 1116
rect 64344 1062 64390 1114
rect 64390 1062 64400 1114
rect 64424 1062 64454 1114
rect 64454 1062 64466 1114
rect 64466 1062 64480 1114
rect 64504 1062 64518 1114
rect 64518 1062 64530 1114
rect 64530 1062 64560 1114
rect 64584 1062 64594 1114
rect 64594 1062 64640 1114
rect 64344 1060 64400 1062
rect 64424 1060 64480 1062
rect 64504 1060 64560 1062
rect 64584 1060 64640 1062
rect 65264 570 65320 572
rect 65344 570 65400 572
rect 65424 570 65480 572
rect 65504 570 65560 572
rect 65264 518 65310 570
rect 65310 518 65320 570
rect 65344 518 65374 570
rect 65374 518 65386 570
rect 65386 518 65400 570
rect 65424 518 65438 570
rect 65438 518 65450 570
rect 65450 518 65480 570
rect 65504 518 65514 570
rect 65514 518 65560 570
rect 65264 516 65320 518
rect 65344 516 65400 518
rect 65424 516 65480 518
rect 65504 516 65560 518
<< metal3 >>
rect 34605 45114 34671 45117
rect 26006 45112 34671 45114
rect 26006 45056 34610 45112
rect 34666 45056 34671 45112
rect 26006 45054 34671 45056
rect 26006 44980 26066 45054
rect 34605 45051 34671 45054
rect 25998 44916 26004 44980
rect 26068 44916 26074 44980
rect 11697 44842 11763 44845
rect 13813 44844 13879 44845
rect 13302 44842 13308 44844
rect 11697 44840 13308 44842
rect 11697 44784 11702 44840
rect 11758 44784 13308 44840
rect 11697 44782 13308 44784
rect 11697 44779 11763 44782
rect 13302 44780 13308 44782
rect 13372 44780 13378 44844
rect 13813 44840 13860 44844
rect 13924 44842 13930 44844
rect 13813 44784 13818 44840
rect 13813 44780 13860 44784
rect 13924 44782 13970 44842
rect 13924 44780 13930 44782
rect 27654 44780 27660 44844
rect 27724 44842 27730 44844
rect 27981 44842 28047 44845
rect 27724 44840 28047 44842
rect 27724 44784 27986 44840
rect 28042 44784 28047 44840
rect 27724 44782 28047 44784
rect 27724 44780 27730 44782
rect 13813 44779 13879 44780
rect 27981 44779 28047 44782
rect 11145 44706 11211 44709
rect 11646 44706 11652 44708
rect 11145 44704 11652 44706
rect 11145 44648 11150 44704
rect 11206 44648 11652 44704
rect 11145 44646 11652 44648
rect 11145 44643 11211 44646
rect 11646 44644 11652 44646
rect 11716 44644 11722 44708
rect 14365 44706 14431 44709
rect 14958 44706 14964 44708
rect 14365 44704 14964 44706
rect 14365 44648 14370 44704
rect 14426 44648 14964 44704
rect 14365 44646 14964 44648
rect 14365 44643 14431 44646
rect 14958 44644 14964 44646
rect 15028 44644 15034 44708
rect 27102 44644 27108 44708
rect 27172 44706 27178 44708
rect 27337 44706 27403 44709
rect 27172 44704 27403 44706
rect 27172 44648 27342 44704
rect 27398 44648 27403 44704
rect 27172 44646 27403 44648
rect 27172 44644 27178 44646
rect 27337 44643 27403 44646
rect 28206 44644 28212 44708
rect 28276 44706 28282 44708
rect 28717 44706 28783 44709
rect 28276 44704 28783 44706
rect 28276 44648 28722 44704
rect 28778 44648 28783 44704
rect 28276 44646 28783 44648
rect 28276 44644 28282 44646
rect 28717 44643 28783 44646
rect 1994 44640 2310 44641
rect 1994 44576 2000 44640
rect 2064 44576 2080 44640
rect 2144 44576 2160 44640
rect 2224 44576 2240 44640
rect 2304 44576 2310 44640
rect 1994 44575 2310 44576
rect 49994 44640 50310 44641
rect 49994 44576 50000 44640
rect 50064 44576 50080 44640
rect 50144 44576 50160 44640
rect 50224 44576 50240 44640
rect 50304 44576 50310 44640
rect 49994 44575 50310 44576
rect 6177 44572 6243 44573
rect 6729 44572 6795 44573
rect 7281 44572 7347 44573
rect 7833 44572 7899 44573
rect 8385 44572 8451 44573
rect 8937 44572 9003 44573
rect 9489 44572 9555 44573
rect 10041 44572 10107 44573
rect 6126 44508 6132 44572
rect 6196 44570 6243 44572
rect 6196 44568 6288 44570
rect 6238 44512 6288 44568
rect 6196 44510 6288 44512
rect 6196 44508 6243 44510
rect 6678 44508 6684 44572
rect 6748 44570 6795 44572
rect 6748 44568 6840 44570
rect 6790 44512 6840 44568
rect 6748 44510 6840 44512
rect 6748 44508 6795 44510
rect 7230 44508 7236 44572
rect 7300 44570 7347 44572
rect 7300 44568 7392 44570
rect 7342 44512 7392 44568
rect 7300 44510 7392 44512
rect 7300 44508 7347 44510
rect 7782 44508 7788 44572
rect 7852 44570 7899 44572
rect 7852 44568 7944 44570
rect 7894 44512 7944 44568
rect 7852 44510 7944 44512
rect 7852 44508 7899 44510
rect 8334 44508 8340 44572
rect 8404 44570 8451 44572
rect 8404 44568 8496 44570
rect 8446 44512 8496 44568
rect 8404 44510 8496 44512
rect 8404 44508 8451 44510
rect 8886 44508 8892 44572
rect 8956 44570 9003 44572
rect 8956 44568 9048 44570
rect 8998 44512 9048 44568
rect 8956 44510 9048 44512
rect 8956 44508 9003 44510
rect 9438 44508 9444 44572
rect 9508 44570 9555 44572
rect 9508 44568 9600 44570
rect 9550 44512 9600 44568
rect 9508 44510 9600 44512
rect 9508 44508 9555 44510
rect 9990 44508 9996 44572
rect 10060 44570 10107 44572
rect 10501 44572 10567 44573
rect 10501 44570 10548 44572
rect 10060 44568 10152 44570
rect 10102 44512 10152 44568
rect 10060 44510 10152 44512
rect 10456 44568 10548 44570
rect 10456 44512 10506 44568
rect 10456 44510 10548 44512
rect 10060 44508 10107 44510
rect 6177 44507 6243 44508
rect 6729 44507 6795 44508
rect 7281 44507 7347 44508
rect 7833 44507 7899 44508
rect 8385 44507 8451 44508
rect 8937 44507 9003 44508
rect 9489 44507 9555 44508
rect 10041 44507 10107 44508
rect 10501 44508 10548 44510
rect 10612 44508 10618 44572
rect 10777 44570 10843 44573
rect 11094 44570 11100 44572
rect 10777 44568 11100 44570
rect 10777 44512 10782 44568
rect 10838 44512 11100 44568
rect 10777 44510 11100 44512
rect 10501 44507 10567 44508
rect 10777 44507 10843 44510
rect 11094 44508 11100 44510
rect 11164 44508 11170 44572
rect 11421 44570 11487 44573
rect 12198 44570 12204 44572
rect 11421 44568 12204 44570
rect 11421 44512 11426 44568
rect 11482 44512 12204 44568
rect 11421 44510 12204 44512
rect 11421 44507 11487 44510
rect 12198 44508 12204 44510
rect 12268 44508 12274 44572
rect 12525 44570 12591 44573
rect 14406 44570 14412 44572
rect 12525 44568 14412 44570
rect 12525 44512 12530 44568
rect 12586 44512 14412 44568
rect 12525 44510 14412 44512
rect 12525 44507 12591 44510
rect 14406 44508 14412 44510
rect 14476 44508 14482 44572
rect 15193 44570 15259 44573
rect 15510 44570 15516 44572
rect 15193 44568 15516 44570
rect 15193 44512 15198 44568
rect 15254 44512 15516 44568
rect 15193 44510 15516 44512
rect 15193 44507 15259 44510
rect 15510 44508 15516 44510
rect 15580 44508 15586 44572
rect 17718 44508 17724 44572
rect 17788 44570 17794 44572
rect 20069 44570 20135 44573
rect 17788 44568 20135 44570
rect 17788 44512 20074 44568
rect 20130 44512 20135 44568
rect 17788 44510 20135 44512
rect 17788 44508 17794 44510
rect 20069 44507 20135 44510
rect 25681 44434 25747 44437
rect 26550 44434 26556 44436
rect 25681 44432 26556 44434
rect 25681 44376 25686 44432
rect 25742 44376 26556 44432
rect 25681 44374 26556 44376
rect 25681 44371 25747 44374
rect 26550 44372 26556 44374
rect 26620 44372 26626 44436
rect 2914 44096 3230 44097
rect 2914 44032 2920 44096
rect 2984 44032 3000 44096
rect 3064 44032 3080 44096
rect 3144 44032 3160 44096
rect 3224 44032 3230 44096
rect 2914 44031 3230 44032
rect 50914 44096 51230 44097
rect 50914 44032 50920 44096
rect 50984 44032 51000 44096
rect 51064 44032 51080 44096
rect 51144 44032 51160 44096
rect 51224 44032 51230 44096
rect 50914 44031 51230 44032
rect 18321 44028 18387 44029
rect 18270 43964 18276 44028
rect 18340 44026 18387 44028
rect 18340 44024 18432 44026
rect 18382 43968 18432 44024
rect 18340 43966 18432 43968
rect 18340 43964 18387 43966
rect 18321 43963 18387 43964
rect 12801 43892 12867 43893
rect 12750 43828 12756 43892
rect 12820 43890 12867 43892
rect 12820 43888 12912 43890
rect 12862 43832 12912 43888
rect 12820 43830 12912 43832
rect 12820 43828 12867 43830
rect 16062 43828 16068 43892
rect 16132 43890 16138 43892
rect 16205 43890 16271 43893
rect 16132 43888 16271 43890
rect 16132 43832 16210 43888
rect 16266 43832 16271 43888
rect 16132 43830 16271 43832
rect 16132 43828 16138 43830
rect 12801 43827 12867 43828
rect 16205 43827 16271 43830
rect 25957 43618 26023 43621
rect 25957 43616 31770 43618
rect 25957 43560 25962 43616
rect 26018 43560 31770 43616
rect 25957 43558 31770 43560
rect 25957 43555 26023 43558
rect 1994 43552 2310 43553
rect 1994 43488 2000 43552
rect 2064 43488 2080 43552
rect 2144 43488 2160 43552
rect 2224 43488 2240 43552
rect 2304 43488 2310 43552
rect 1994 43487 2310 43488
rect 17166 43420 17172 43484
rect 17236 43482 17242 43484
rect 17493 43482 17559 43485
rect 17236 43480 17559 43482
rect 17236 43424 17498 43480
rect 17554 43424 17559 43480
rect 17236 43422 17559 43424
rect 17236 43420 17242 43422
rect 17493 43419 17559 43422
rect 23238 43420 23244 43484
rect 23308 43482 23314 43484
rect 31710 43482 31770 43558
rect 49994 43552 50310 43553
rect 49994 43488 50000 43552
rect 50064 43488 50080 43552
rect 50144 43488 50160 43552
rect 50224 43488 50240 43552
rect 50304 43488 50310 43552
rect 49994 43487 50310 43488
rect 32070 43482 32076 43484
rect 23308 43422 26250 43482
rect 31710 43422 32076 43482
rect 23308 43420 23314 43422
rect 22134 43284 22140 43348
rect 22204 43346 22210 43348
rect 24710 43346 24716 43348
rect 22204 43286 24716 43346
rect 22204 43284 22210 43286
rect 24710 43284 24716 43286
rect 24780 43284 24786 43348
rect 26190 43346 26250 43422
rect 32070 43420 32076 43422
rect 32140 43420 32146 43484
rect 34237 43346 34303 43349
rect 26190 43344 34303 43346
rect 26190 43288 34242 43344
rect 34298 43288 34303 43344
rect 26190 43286 34303 43288
rect 34237 43283 34303 43286
rect 20437 43210 20503 43213
rect 35198 43210 35204 43212
rect 20437 43208 35204 43210
rect 20437 43152 20442 43208
rect 20498 43152 35204 43208
rect 20437 43150 35204 43152
rect 20437 43147 20503 43150
rect 35198 43148 35204 43150
rect 35268 43148 35274 43212
rect 24945 43074 25011 43077
rect 25497 43074 25563 43077
rect 27470 43074 27476 43076
rect 24945 43072 27476 43074
rect 24945 43016 24950 43072
rect 25006 43016 25502 43072
rect 25558 43016 27476 43072
rect 24945 43014 27476 43016
rect 24945 43011 25011 43014
rect 25497 43011 25563 43014
rect 27470 43012 27476 43014
rect 27540 43012 27546 43076
rect 27654 43012 27660 43076
rect 27724 43074 27730 43076
rect 36169 43074 36235 43077
rect 27724 43072 36235 43074
rect 27724 43016 36174 43072
rect 36230 43016 36235 43072
rect 27724 43014 36235 43016
rect 27724 43012 27730 43014
rect 36169 43011 36235 43014
rect 41781 43074 41847 43077
rect 44265 43074 44331 43077
rect 41781 43072 44331 43074
rect 41781 43016 41786 43072
rect 41842 43016 44270 43072
rect 44326 43016 44331 43072
rect 41781 43014 44331 43016
rect 41781 43011 41847 43014
rect 44265 43011 44331 43014
rect 2914 43008 3230 43009
rect 2914 42944 2920 43008
rect 2984 42944 3000 43008
rect 3064 42944 3080 43008
rect 3144 42944 3160 43008
rect 3224 42944 3230 43008
rect 2914 42943 3230 42944
rect 50914 43008 51230 43009
rect 50914 42944 50920 43008
rect 50984 42944 51000 43008
rect 51064 42944 51080 43008
rect 51144 42944 51160 43008
rect 51224 42944 51230 43008
rect 50914 42943 51230 42944
rect 16614 42876 16620 42940
rect 16684 42938 16690 42940
rect 17309 42938 17375 42941
rect 16684 42936 17375 42938
rect 16684 42880 17314 42936
rect 17370 42880 17375 42936
rect 16684 42878 17375 42880
rect 16684 42876 16690 42878
rect 17309 42875 17375 42878
rect 24894 42876 24900 42940
rect 24964 42938 24970 42940
rect 26141 42938 26207 42941
rect 24964 42936 26207 42938
rect 24964 42880 26146 42936
rect 26202 42880 26207 42936
rect 24964 42878 26207 42880
rect 24964 42876 24970 42878
rect 26141 42875 26207 42878
rect 21357 42666 21423 42669
rect 24209 42666 24275 42669
rect 21357 42664 24275 42666
rect 21357 42608 21362 42664
rect 21418 42608 24214 42664
rect 24270 42608 24275 42664
rect 21357 42606 24275 42608
rect 21357 42603 21423 42606
rect 24209 42603 24275 42606
rect 25313 42666 25379 42669
rect 47393 42666 47459 42669
rect 25313 42664 47459 42666
rect 25313 42608 25318 42664
rect 25374 42608 47398 42664
rect 47454 42608 47459 42664
rect 25313 42606 47459 42608
rect 25313 42603 25379 42606
rect 47393 42603 47459 42606
rect 1994 42464 2310 42465
rect 1994 42400 2000 42464
rect 2064 42400 2080 42464
rect 2144 42400 2160 42464
rect 2224 42400 2240 42464
rect 2304 42400 2310 42464
rect 1994 42399 2310 42400
rect 49994 42464 50310 42465
rect 49994 42400 50000 42464
rect 50064 42400 50080 42464
rect 50144 42400 50160 42464
rect 50224 42400 50240 42464
rect 50304 42400 50310 42464
rect 49994 42399 50310 42400
rect 17953 42394 18019 42397
rect 18822 42394 18828 42396
rect 17953 42392 18828 42394
rect 17953 42336 17958 42392
rect 18014 42336 18828 42392
rect 17953 42334 18828 42336
rect 17953 42331 18019 42334
rect 18822 42332 18828 42334
rect 18892 42332 18898 42396
rect 37089 42394 37155 42397
rect 22050 42392 37155 42394
rect 22050 42336 37094 42392
rect 37150 42336 37155 42392
rect 22050 42334 37155 42336
rect 15561 42258 15627 42261
rect 22050 42258 22110 42334
rect 37089 42331 37155 42334
rect 15561 42256 22110 42258
rect 15561 42200 15566 42256
rect 15622 42200 22110 42256
rect 15561 42198 22110 42200
rect 35893 42258 35959 42261
rect 58065 42258 58131 42261
rect 35893 42256 58131 42258
rect 35893 42200 35898 42256
rect 35954 42200 58070 42256
rect 58126 42200 58131 42256
rect 35893 42198 58131 42200
rect 15561 42195 15627 42198
rect 35893 42195 35959 42198
rect 58065 42195 58131 42198
rect 17953 42122 18019 42125
rect 30649 42122 30715 42125
rect 30966 42122 30972 42124
rect 17953 42120 29930 42122
rect 17953 42064 17958 42120
rect 18014 42064 29930 42120
rect 17953 42062 29930 42064
rect 17953 42059 18019 42062
rect 25221 41986 25287 41989
rect 29637 41986 29703 41989
rect 25221 41984 29703 41986
rect 25221 41928 25226 41984
rect 25282 41928 29642 41984
rect 29698 41928 29703 41984
rect 25221 41926 29703 41928
rect 29870 41986 29930 42062
rect 30649 42120 30972 42122
rect 30649 42064 30654 42120
rect 30710 42064 30972 42120
rect 30649 42062 30972 42064
rect 30649 42059 30715 42062
rect 30966 42060 30972 42062
rect 31036 42060 31042 42124
rect 32029 42122 32095 42125
rect 44265 42122 44331 42125
rect 32029 42120 44331 42122
rect 32029 42064 32034 42120
rect 32090 42064 44270 42120
rect 44326 42064 44331 42120
rect 32029 42062 44331 42064
rect 32029 42059 32095 42062
rect 44265 42059 44331 42062
rect 30649 41986 30715 41989
rect 29870 41984 30715 41986
rect 29870 41928 30654 41984
rect 30710 41928 30715 41984
rect 29870 41926 30715 41928
rect 25221 41923 25287 41926
rect 29637 41923 29703 41926
rect 30649 41923 30715 41926
rect 2914 41920 3230 41921
rect 2914 41856 2920 41920
rect 2984 41856 3000 41920
rect 3064 41856 3080 41920
rect 3144 41856 3160 41920
rect 3224 41856 3230 41920
rect 2914 41855 3230 41856
rect 50914 41920 51230 41921
rect 50914 41856 50920 41920
rect 50984 41856 51000 41920
rect 51064 41856 51080 41920
rect 51144 41856 51160 41920
rect 51224 41856 51230 41920
rect 50914 41855 51230 41856
rect 25497 41850 25563 41853
rect 43069 41850 43135 41853
rect 25497 41848 43135 41850
rect 25497 41792 25502 41848
rect 25558 41792 43074 41848
rect 43130 41792 43135 41848
rect 25497 41790 43135 41792
rect 25497 41787 25563 41790
rect 43069 41787 43135 41790
rect 22093 41714 22159 41717
rect 22369 41714 22435 41717
rect 22093 41712 22435 41714
rect 22093 41656 22098 41712
rect 22154 41656 22374 41712
rect 22430 41656 22435 41712
rect 22093 41654 22435 41656
rect 22093 41651 22159 41654
rect 22369 41651 22435 41654
rect 23105 41714 23171 41717
rect 25773 41714 25839 41717
rect 23105 41712 25839 41714
rect 23105 41656 23110 41712
rect 23166 41656 25778 41712
rect 25834 41656 25839 41712
rect 23105 41654 25839 41656
rect 23105 41651 23171 41654
rect 25773 41651 25839 41654
rect 26049 41714 26115 41717
rect 29177 41714 29243 41717
rect 26049 41712 29243 41714
rect 26049 41656 26054 41712
rect 26110 41656 29182 41712
rect 29238 41656 29243 41712
rect 26049 41654 29243 41656
rect 26049 41651 26115 41654
rect 29177 41651 29243 41654
rect 30373 41714 30439 41717
rect 43529 41714 43595 41717
rect 30373 41712 43595 41714
rect 30373 41656 30378 41712
rect 30434 41656 43534 41712
rect 43590 41656 43595 41712
rect 30373 41654 43595 41656
rect 30373 41651 30439 41654
rect 43529 41651 43595 41654
rect 24669 41578 24735 41581
rect 30373 41578 30439 41581
rect 60733 41578 60799 41581
rect 24669 41576 26618 41578
rect 24669 41520 24674 41576
rect 24730 41520 26618 41576
rect 24669 41518 26618 41520
rect 24669 41515 24735 41518
rect 26049 41442 26115 41445
rect 26558 41442 26618 41518
rect 30373 41576 60799 41578
rect 30373 41520 30378 41576
rect 30434 41520 60738 41576
rect 60794 41520 60799 41576
rect 30373 41518 60799 41520
rect 30373 41515 30439 41518
rect 60733 41515 60799 41518
rect 34789 41442 34855 41445
rect 26049 41440 26434 41442
rect 26049 41384 26054 41440
rect 26110 41384 26434 41440
rect 26049 41382 26434 41384
rect 26558 41440 34855 41442
rect 26558 41384 34794 41440
rect 34850 41384 34855 41440
rect 26558 41382 34855 41384
rect 26049 41379 26115 41382
rect 1994 41376 2310 41377
rect 1994 41312 2000 41376
rect 2064 41312 2080 41376
rect 2144 41312 2160 41376
rect 2224 41312 2240 41376
rect 2304 41312 2310 41376
rect 1994 41311 2310 41312
rect 25865 41306 25931 41309
rect 26374 41306 26434 41382
rect 34789 41379 34855 41382
rect 49994 41376 50310 41377
rect 49994 41312 50000 41376
rect 50064 41312 50080 41376
rect 50144 41312 50160 41376
rect 50224 41312 50240 41376
rect 50304 41312 50310 41376
rect 49994 41311 50310 41312
rect 25865 41304 26434 41306
rect 25865 41248 25870 41304
rect 25926 41248 26434 41304
rect 25865 41246 26434 41248
rect 30649 41306 30715 41309
rect 35014 41306 35020 41308
rect 30649 41304 35020 41306
rect 30649 41248 30654 41304
rect 30710 41248 35020 41304
rect 30649 41246 35020 41248
rect 25865 41243 25931 41246
rect 30649 41243 30715 41246
rect 35014 41244 35020 41246
rect 35084 41244 35090 41308
rect 40677 41306 40743 41309
rect 43897 41306 43963 41309
rect 40677 41304 43963 41306
rect 40677 41248 40682 41304
rect 40738 41248 43902 41304
rect 43958 41248 43963 41304
rect 40677 41246 43963 41248
rect 40677 41243 40743 41246
rect 43897 41243 43963 41246
rect 30373 41170 30439 41173
rect 26558 41168 30439 41170
rect 26558 41112 30378 41168
rect 30434 41112 30439 41168
rect 26558 41110 30439 41112
rect 13997 41034 14063 41037
rect 25957 41034 26023 41037
rect 13997 41032 26023 41034
rect 13997 40976 14002 41032
rect 14058 40976 25962 41032
rect 26018 40976 26023 41032
rect 13997 40974 26023 40976
rect 13997 40971 14063 40974
rect 25957 40971 26023 40974
rect 26141 41034 26207 41037
rect 26558 41034 26618 41110
rect 30373 41107 30439 41110
rect 33317 41170 33383 41173
rect 63585 41170 63651 41173
rect 33317 41168 63651 41170
rect 33317 41112 33322 41168
rect 33378 41112 63590 41168
rect 63646 41112 63651 41168
rect 33317 41110 63651 41112
rect 33317 41107 33383 41110
rect 63585 41107 63651 41110
rect 26141 41032 26618 41034
rect 26141 40976 26146 41032
rect 26202 40976 26618 41032
rect 26141 40974 26618 40976
rect 26141 40971 26207 40974
rect 26918 40972 26924 41036
rect 26988 41034 26994 41036
rect 36721 41034 36787 41037
rect 26988 41032 36787 41034
rect 26988 40976 36726 41032
rect 36782 40976 36787 41032
rect 26988 40974 36787 40976
rect 26988 40972 26994 40974
rect 36721 40971 36787 40974
rect 50889 41034 50955 41037
rect 55765 41034 55831 41037
rect 56593 41034 56659 41037
rect 50889 41032 56659 41034
rect 50889 40976 50894 41032
rect 50950 40976 55770 41032
rect 55826 40976 56598 41032
rect 56654 40976 56659 41032
rect 50889 40974 56659 40976
rect 50889 40971 50955 40974
rect 55765 40971 55831 40974
rect 56593 40971 56659 40974
rect 22645 40898 22711 40901
rect 32990 40898 32996 40900
rect 22645 40896 32996 40898
rect 22645 40840 22650 40896
rect 22706 40840 32996 40896
rect 22645 40838 32996 40840
rect 22645 40835 22711 40838
rect 32990 40836 32996 40838
rect 33060 40836 33066 40900
rect 2914 40832 3230 40833
rect 2914 40768 2920 40832
rect 2984 40768 3000 40832
rect 3064 40768 3080 40832
rect 3144 40768 3160 40832
rect 3224 40768 3230 40832
rect 2914 40767 3230 40768
rect 50914 40832 51230 40833
rect 50914 40768 50920 40832
rect 50984 40768 51000 40832
rect 51064 40768 51080 40832
rect 51144 40768 51160 40832
rect 51224 40768 51230 40832
rect 50914 40767 51230 40768
rect 27470 40700 27476 40764
rect 27540 40762 27546 40764
rect 41965 40762 42031 40765
rect 27540 40760 42031 40762
rect 27540 40704 41970 40760
rect 42026 40704 42031 40760
rect 27540 40702 42031 40704
rect 27540 40700 27546 40702
rect 41965 40699 42031 40702
rect 3918 40564 3924 40628
rect 3988 40626 3994 40628
rect 23790 40626 23796 40628
rect 3988 40566 23796 40626
rect 3988 40564 3994 40566
rect 23790 40564 23796 40566
rect 23860 40564 23866 40628
rect 25446 40564 25452 40628
rect 25516 40626 25522 40628
rect 32806 40626 32812 40628
rect 25516 40566 32812 40626
rect 25516 40564 25522 40566
rect 32806 40564 32812 40566
rect 32876 40564 32882 40628
rect 34421 40626 34487 40629
rect 47853 40626 47919 40629
rect 48221 40626 48287 40629
rect 34421 40624 48287 40626
rect 34421 40568 34426 40624
rect 34482 40568 47858 40624
rect 47914 40568 48226 40624
rect 48282 40568 48287 40624
rect 34421 40566 48287 40568
rect 34421 40563 34487 40566
rect 47853 40563 47919 40566
rect 48221 40563 48287 40566
rect 20805 40490 20871 40493
rect 49785 40490 49851 40493
rect 20805 40488 49851 40490
rect 20805 40432 20810 40488
rect 20866 40432 49790 40488
rect 49846 40432 49851 40488
rect 20805 40430 49851 40432
rect 20805 40427 20871 40430
rect 49785 40427 49851 40430
rect 18505 40354 18571 40357
rect 27838 40354 27844 40356
rect 18505 40352 27844 40354
rect 18505 40296 18510 40352
rect 18566 40296 27844 40352
rect 18505 40294 27844 40296
rect 18505 40291 18571 40294
rect 27838 40292 27844 40294
rect 27908 40292 27914 40356
rect 1994 40288 2310 40289
rect 1994 40224 2000 40288
rect 2064 40224 2080 40288
rect 2144 40224 2160 40288
rect 2224 40224 2240 40288
rect 2304 40224 2310 40288
rect 1994 40223 2310 40224
rect 49994 40288 50310 40289
rect 49994 40224 50000 40288
rect 50064 40224 50080 40288
rect 50144 40224 50160 40288
rect 50224 40224 50240 40288
rect 50304 40224 50310 40288
rect 49994 40223 50310 40224
rect 31293 40218 31359 40221
rect 38837 40218 38903 40221
rect 27662 40216 31359 40218
rect 27662 40160 31298 40216
rect 31354 40160 31359 40216
rect 27662 40158 31359 40160
rect 24342 40020 24348 40084
rect 24412 40082 24418 40084
rect 25037 40082 25103 40085
rect 24412 40080 25103 40082
rect 24412 40024 25042 40080
rect 25098 40024 25103 40080
rect 24412 40022 25103 40024
rect 24412 40020 24418 40022
rect 25037 40019 25103 40022
rect 13629 39946 13695 39949
rect 27662 39946 27722 40158
rect 31293 40155 31359 40158
rect 31710 40216 38903 40218
rect 31710 40160 38842 40216
rect 38898 40160 38903 40216
rect 31710 40158 38903 40160
rect 31710 40082 31770 40158
rect 38837 40155 38903 40158
rect 30284 40022 31770 40082
rect 34697 40082 34763 40085
rect 62665 40082 62731 40085
rect 34697 40080 62731 40082
rect 34697 40024 34702 40080
rect 34758 40024 62670 40080
rect 62726 40024 62731 40080
rect 34697 40022 62731 40024
rect 13629 39944 27722 39946
rect 13629 39888 13634 39944
rect 13690 39888 27722 39944
rect 13629 39886 27722 39888
rect 13629 39883 13695 39886
rect 28574 39884 28580 39948
rect 28644 39946 28650 39948
rect 30284 39946 30344 40022
rect 34697 40019 34763 40022
rect 62665 40019 62731 40022
rect 28644 39886 30344 39946
rect 31845 39946 31911 39949
rect 35801 39946 35867 39949
rect 31845 39944 35867 39946
rect 31845 39888 31850 39944
rect 31906 39888 35806 39944
rect 35862 39888 35867 39944
rect 31845 39886 35867 39888
rect 28644 39884 28650 39886
rect 31845 39883 31911 39886
rect 35801 39883 35867 39886
rect 15510 39748 15516 39812
rect 15580 39810 15586 39812
rect 34421 39810 34487 39813
rect 15580 39808 34487 39810
rect 15580 39752 34426 39808
rect 34482 39752 34487 39808
rect 15580 39750 34487 39752
rect 15580 39748 15586 39750
rect 34421 39747 34487 39750
rect 41045 39810 41111 39813
rect 44725 39810 44791 39813
rect 41045 39808 44791 39810
rect 41045 39752 41050 39808
rect 41106 39752 44730 39808
rect 44786 39752 44791 39808
rect 41045 39750 44791 39752
rect 41045 39747 41111 39750
rect 44725 39747 44791 39750
rect 2914 39744 3230 39745
rect 2914 39680 2920 39744
rect 2984 39680 3000 39744
rect 3064 39680 3080 39744
rect 3144 39680 3160 39744
rect 3224 39680 3230 39744
rect 2914 39679 3230 39680
rect 50914 39744 51230 39745
rect 50914 39680 50920 39744
rect 50984 39680 51000 39744
rect 51064 39680 51080 39744
rect 51144 39680 51160 39744
rect 51224 39680 51230 39744
rect 50914 39679 51230 39680
rect 11421 39674 11487 39677
rect 27613 39674 27679 39677
rect 11421 39672 27679 39674
rect 11421 39616 11426 39672
rect 11482 39616 27618 39672
rect 27674 39616 27679 39672
rect 11421 39614 27679 39616
rect 11421 39611 11487 39614
rect 27613 39611 27679 39614
rect 32990 39612 32996 39676
rect 33060 39674 33066 39676
rect 36118 39674 36124 39676
rect 33060 39614 36124 39674
rect 33060 39612 33066 39614
rect 36118 39612 36124 39614
rect 36188 39612 36194 39676
rect 36629 39674 36695 39677
rect 38745 39674 38811 39677
rect 36629 39672 38811 39674
rect 36629 39616 36634 39672
rect 36690 39616 38750 39672
rect 38806 39616 38811 39672
rect 36629 39614 38811 39616
rect 36629 39611 36695 39614
rect 38745 39611 38811 39614
rect 25037 39538 25103 39541
rect 52545 39538 52611 39541
rect 52821 39538 52887 39541
rect 25037 39536 52887 39538
rect 25037 39480 25042 39536
rect 25098 39480 52550 39536
rect 52606 39480 52826 39536
rect 52882 39480 52887 39536
rect 25037 39478 52887 39480
rect 25037 39475 25103 39478
rect 52545 39475 52611 39478
rect 52821 39475 52887 39478
rect 19006 39340 19012 39404
rect 19076 39402 19082 39404
rect 45093 39402 45159 39405
rect 64689 39402 64755 39405
rect 19076 39400 45159 39402
rect 19076 39344 45098 39400
rect 45154 39344 45159 39400
rect 19076 39342 45159 39344
rect 19076 39340 19082 39342
rect 45093 39339 45159 39342
rect 46246 39400 64755 39402
rect 46246 39344 64694 39400
rect 64750 39344 64755 39400
rect 46246 39342 64755 39344
rect 21173 39266 21239 39269
rect 25037 39266 25103 39269
rect 21173 39264 25103 39266
rect 21173 39208 21178 39264
rect 21234 39208 25042 39264
rect 25098 39208 25103 39264
rect 21173 39206 25103 39208
rect 21173 39203 21239 39206
rect 25037 39203 25103 39206
rect 27838 39204 27844 39268
rect 27908 39266 27914 39268
rect 31569 39266 31635 39269
rect 27908 39264 31635 39266
rect 27908 39208 31574 39264
rect 31630 39208 31635 39264
rect 27908 39206 31635 39208
rect 27908 39204 27914 39206
rect 31569 39203 31635 39206
rect 32806 39204 32812 39268
rect 32876 39266 32882 39268
rect 36721 39266 36787 39269
rect 32876 39264 36787 39266
rect 32876 39208 36726 39264
rect 36782 39208 36787 39264
rect 32876 39206 36787 39208
rect 32876 39204 32882 39206
rect 36721 39203 36787 39206
rect 41229 39266 41295 39269
rect 41597 39266 41663 39269
rect 41229 39264 41663 39266
rect 41229 39208 41234 39264
rect 41290 39208 41602 39264
rect 41658 39208 41663 39264
rect 41229 39206 41663 39208
rect 41229 39203 41295 39206
rect 41597 39203 41663 39206
rect 1994 39200 2310 39201
rect 1994 39136 2000 39200
rect 2064 39136 2080 39200
rect 2144 39136 2160 39200
rect 2224 39136 2240 39200
rect 2304 39136 2310 39200
rect 1994 39135 2310 39136
rect 30373 39130 30439 39133
rect 46246 39130 46306 39342
rect 64689 39339 64755 39342
rect 49994 39200 50310 39201
rect 49994 39136 50000 39200
rect 50064 39136 50080 39200
rect 50144 39136 50160 39200
rect 50224 39136 50240 39200
rect 50304 39136 50310 39200
rect 49994 39135 50310 39136
rect 30373 39128 46306 39130
rect 30373 39072 30378 39128
rect 30434 39072 46306 39128
rect 30373 39070 46306 39072
rect 30373 39067 30439 39070
rect 21081 38994 21147 38997
rect 27981 38994 28047 38997
rect 21081 38992 28047 38994
rect 21081 38936 21086 38992
rect 21142 38936 27986 38992
rect 28042 38936 28047 38992
rect 21081 38934 28047 38936
rect 21081 38931 21147 38934
rect 27981 38931 28047 38934
rect 28942 38932 28948 38996
rect 29012 38994 29018 38996
rect 31385 38994 31451 38997
rect 29012 38992 31451 38994
rect 29012 38936 31390 38992
rect 31446 38936 31451 38992
rect 29012 38934 31451 38936
rect 29012 38932 29018 38934
rect 31385 38931 31451 38934
rect 33041 38994 33107 38997
rect 33041 38992 60750 38994
rect 33041 38936 33046 38992
rect 33102 38936 60750 38992
rect 33041 38934 60750 38936
rect 33041 38931 33107 38934
rect 16205 38858 16271 38861
rect 52085 38858 52151 38861
rect 16205 38856 52151 38858
rect 16205 38800 16210 38856
rect 16266 38800 52090 38856
rect 52146 38800 52151 38856
rect 16205 38798 52151 38800
rect 16205 38795 16271 38798
rect 52085 38795 52151 38798
rect 26182 38660 26188 38724
rect 26252 38722 26258 38724
rect 26601 38722 26667 38725
rect 26252 38720 26667 38722
rect 26252 38664 26606 38720
rect 26662 38664 26667 38720
rect 26252 38662 26667 38664
rect 26252 38660 26258 38662
rect 26601 38659 26667 38662
rect 28390 38660 28396 38724
rect 28460 38722 28466 38724
rect 31937 38722 32003 38725
rect 28460 38720 32003 38722
rect 28460 38664 31942 38720
rect 31998 38664 32003 38720
rect 28460 38662 32003 38664
rect 28460 38660 28466 38662
rect 31937 38659 32003 38662
rect 32121 38722 32187 38725
rect 32438 38722 32444 38724
rect 32121 38720 32444 38722
rect 32121 38664 32126 38720
rect 32182 38664 32444 38720
rect 32121 38662 32444 38664
rect 32121 38659 32187 38662
rect 32438 38660 32444 38662
rect 32508 38660 32514 38724
rect 33174 38722 33180 38724
rect 32878 38662 33180 38722
rect 2914 38656 3230 38657
rect 2914 38592 2920 38656
rect 2984 38592 3000 38656
rect 3064 38592 3080 38656
rect 3144 38592 3160 38656
rect 3224 38592 3230 38656
rect 2914 38591 3230 38592
rect 24577 38588 24643 38589
rect 24526 38586 24532 38588
rect 24486 38526 24532 38586
rect 24596 38584 24643 38588
rect 24638 38528 24643 38584
rect 24526 38524 24532 38526
rect 24596 38524 24643 38528
rect 24577 38523 24643 38524
rect 27429 38586 27495 38589
rect 30833 38586 30899 38589
rect 32878 38586 32938 38662
rect 33174 38660 33180 38662
rect 33244 38660 33250 38724
rect 33593 38722 33659 38725
rect 35382 38722 35388 38724
rect 33593 38720 35388 38722
rect 33593 38664 33598 38720
rect 33654 38664 35388 38720
rect 33593 38662 35388 38664
rect 33593 38659 33659 38662
rect 35382 38660 35388 38662
rect 35452 38660 35458 38724
rect 43897 38722 43963 38725
rect 46974 38722 46980 38724
rect 43897 38720 46980 38722
rect 43897 38664 43902 38720
rect 43958 38664 46980 38720
rect 43897 38662 46980 38664
rect 43897 38659 43963 38662
rect 46974 38660 46980 38662
rect 47044 38660 47050 38724
rect 50914 38656 51230 38657
rect 50914 38592 50920 38656
rect 50984 38592 51000 38656
rect 51064 38592 51080 38656
rect 51144 38592 51160 38656
rect 51224 38592 51230 38656
rect 50914 38591 51230 38592
rect 34094 38586 34100 38588
rect 27429 38584 30482 38586
rect 27429 38528 27434 38584
rect 27490 38528 30482 38584
rect 27429 38526 30482 38528
rect 27429 38523 27495 38526
rect 25998 38388 26004 38452
rect 26068 38450 26074 38452
rect 28533 38450 28599 38453
rect 26068 38448 28599 38450
rect 26068 38392 28538 38448
rect 28594 38392 28599 38448
rect 26068 38390 28599 38392
rect 30422 38450 30482 38526
rect 30833 38584 32938 38586
rect 30833 38528 30838 38584
rect 30894 38528 32938 38584
rect 30833 38526 32938 38528
rect 33016 38526 34100 38586
rect 30833 38523 30899 38526
rect 33016 38450 33076 38526
rect 34094 38524 34100 38526
rect 34164 38524 34170 38588
rect 34973 38586 35039 38589
rect 35617 38586 35683 38589
rect 34973 38584 35683 38586
rect 34973 38528 34978 38584
rect 35034 38528 35622 38584
rect 35678 38528 35683 38584
rect 34973 38526 35683 38528
rect 34973 38523 35039 38526
rect 35617 38523 35683 38526
rect 41045 38586 41111 38589
rect 45093 38586 45159 38589
rect 41045 38584 45159 38586
rect 41045 38528 41050 38584
rect 41106 38528 45098 38584
rect 45154 38528 45159 38584
rect 41045 38526 45159 38528
rect 41045 38523 41111 38526
rect 45093 38523 45159 38526
rect 48313 38586 48379 38589
rect 48865 38586 48931 38589
rect 49969 38586 50035 38589
rect 48313 38584 50035 38586
rect 48313 38528 48318 38584
rect 48374 38528 48870 38584
rect 48926 38528 49974 38584
rect 50030 38528 50035 38584
rect 48313 38526 50035 38528
rect 60690 38586 60750 38934
rect 62798 38586 62804 38588
rect 60690 38526 62804 38586
rect 48313 38523 48379 38526
rect 48865 38523 48931 38526
rect 49969 38523 50035 38526
rect 62798 38524 62804 38526
rect 62868 38524 62874 38588
rect 30422 38390 33076 38450
rect 33225 38450 33291 38453
rect 55213 38450 55279 38453
rect 33225 38448 55279 38450
rect 33225 38392 33230 38448
rect 33286 38392 55218 38448
rect 55274 38392 55279 38448
rect 33225 38390 55279 38392
rect 26068 38388 26074 38390
rect 28533 38387 28599 38390
rect 33225 38387 33291 38390
rect 55213 38387 55279 38390
rect 21398 38252 21404 38316
rect 21468 38314 21474 38316
rect 41965 38314 42031 38317
rect 21468 38312 42031 38314
rect 21468 38256 41970 38312
rect 42026 38256 42031 38312
rect 21468 38254 42031 38256
rect 21468 38252 21474 38254
rect 41965 38251 42031 38254
rect 26693 38178 26759 38181
rect 28349 38178 28415 38181
rect 26693 38176 28415 38178
rect 26693 38120 26698 38176
rect 26754 38120 28354 38176
rect 28410 38120 28415 38176
rect 26693 38118 28415 38120
rect 26693 38115 26759 38118
rect 28349 38115 28415 38118
rect 28533 38178 28599 38181
rect 33133 38178 33199 38181
rect 28533 38176 33199 38178
rect 28533 38120 28538 38176
rect 28594 38120 33138 38176
rect 33194 38120 33199 38176
rect 28533 38118 33199 38120
rect 28533 38115 28599 38118
rect 33133 38115 33199 38118
rect 33685 38178 33751 38181
rect 33685 38176 46306 38178
rect 33685 38120 33690 38176
rect 33746 38120 46306 38176
rect 33685 38118 46306 38120
rect 33685 38115 33751 38118
rect 1994 38112 2310 38113
rect 1994 38048 2000 38112
rect 2064 38048 2080 38112
rect 2144 38048 2160 38112
rect 2224 38048 2240 38112
rect 2304 38048 2310 38112
rect 1994 38047 2310 38048
rect 20110 37980 20116 38044
rect 20180 38042 20186 38044
rect 44541 38042 44607 38045
rect 20180 38040 44607 38042
rect 20180 37984 44546 38040
rect 44602 37984 44607 38040
rect 20180 37982 44607 37984
rect 20180 37980 20186 37982
rect 44541 37979 44607 37982
rect 16573 37906 16639 37909
rect 27797 37906 27863 37909
rect 16573 37904 27863 37906
rect 16573 37848 16578 37904
rect 16634 37848 27802 37904
rect 27858 37848 27863 37904
rect 16573 37846 27863 37848
rect 16573 37843 16639 37846
rect 27797 37843 27863 37846
rect 28022 37844 28028 37908
rect 28092 37906 28098 37908
rect 30833 37906 30899 37909
rect 28092 37904 30899 37906
rect 28092 37848 30838 37904
rect 30894 37848 30899 37904
rect 28092 37846 30899 37848
rect 28092 37844 28098 37846
rect 30833 37843 30899 37846
rect 31477 37906 31543 37909
rect 34237 37906 34303 37909
rect 31477 37904 34303 37906
rect 31477 37848 31482 37904
rect 31538 37848 34242 37904
rect 34298 37848 34303 37904
rect 31477 37846 34303 37848
rect 31477 37843 31543 37846
rect 34237 37843 34303 37846
rect 39665 37906 39731 37909
rect 41321 37906 41387 37909
rect 39665 37904 41387 37906
rect 39665 37848 39670 37904
rect 39726 37848 41326 37904
rect 41382 37848 41387 37904
rect 39665 37846 41387 37848
rect 46246 37906 46306 38118
rect 49994 38112 50310 38113
rect 49994 38048 50000 38112
rect 50064 38048 50080 38112
rect 50144 38048 50160 38112
rect 50224 38048 50240 38112
rect 50304 38048 50310 38112
rect 49994 38047 50310 38048
rect 56685 37906 56751 37909
rect 46246 37904 56751 37906
rect 46246 37848 56690 37904
rect 56746 37848 56751 37904
rect 46246 37846 56751 37848
rect 39665 37843 39731 37846
rect 41321 37843 41387 37846
rect 56685 37843 56751 37846
rect 18045 37770 18111 37773
rect 26693 37770 26759 37773
rect 28073 37770 28139 37773
rect 18045 37768 26759 37770
rect 18045 37712 18050 37768
rect 18106 37712 26698 37768
rect 26754 37712 26759 37768
rect 18045 37710 26759 37712
rect 18045 37707 18111 37710
rect 26693 37707 26759 37710
rect 26926 37768 28139 37770
rect 26926 37712 28078 37768
rect 28134 37712 28139 37768
rect 26926 37710 28139 37712
rect 17953 37634 18019 37637
rect 26926 37634 26986 37710
rect 28073 37707 28139 37710
rect 28349 37770 28415 37773
rect 33225 37770 33291 37773
rect 33685 37770 33751 37773
rect 28349 37768 33751 37770
rect 28349 37712 28354 37768
rect 28410 37712 33230 37768
rect 33286 37712 33690 37768
rect 33746 37712 33751 37768
rect 28349 37710 33751 37712
rect 28349 37707 28415 37710
rect 33225 37707 33291 37710
rect 33685 37707 33751 37710
rect 34697 37770 34763 37773
rect 62982 37770 62988 37772
rect 34697 37768 62988 37770
rect 34697 37712 34702 37768
rect 34758 37712 62988 37768
rect 34697 37710 62988 37712
rect 34697 37707 34763 37710
rect 62982 37708 62988 37710
rect 63052 37708 63058 37772
rect 17953 37632 26986 37634
rect 17953 37576 17958 37632
rect 18014 37576 26986 37632
rect 17953 37574 26986 37576
rect 27521 37634 27587 37637
rect 35341 37634 35407 37637
rect 27521 37632 35407 37634
rect 27521 37576 27526 37632
rect 27582 37576 35346 37632
rect 35402 37576 35407 37632
rect 27521 37574 35407 37576
rect 17953 37571 18019 37574
rect 27521 37571 27587 37574
rect 35341 37571 35407 37574
rect 2914 37568 3230 37569
rect 2914 37504 2920 37568
rect 2984 37504 3000 37568
rect 3064 37504 3080 37568
rect 3144 37504 3160 37568
rect 3224 37504 3230 37568
rect 2914 37503 3230 37504
rect 50914 37568 51230 37569
rect 50914 37504 50920 37568
rect 50984 37504 51000 37568
rect 51064 37504 51080 37568
rect 51144 37504 51160 37568
rect 51224 37504 51230 37568
rect 50914 37503 51230 37504
rect 65254 37568 65570 37569
rect 65254 37504 65260 37568
rect 65324 37504 65340 37568
rect 65404 37504 65420 37568
rect 65484 37504 65500 37568
rect 65564 37504 65570 37568
rect 65254 37503 65570 37504
rect 12617 37498 12683 37501
rect 25773 37498 25839 37501
rect 12617 37496 25839 37498
rect 12617 37440 12622 37496
rect 12678 37440 25778 37496
rect 25834 37440 25839 37496
rect 12617 37438 25839 37440
rect 12617 37435 12683 37438
rect 25773 37435 25839 37438
rect 27286 37436 27292 37500
rect 27356 37498 27362 37500
rect 28349 37498 28415 37501
rect 27356 37496 28415 37498
rect 27356 37440 28354 37496
rect 28410 37440 28415 37496
rect 27356 37438 28415 37440
rect 27356 37436 27362 37438
rect 28349 37435 28415 37438
rect 28533 37500 28599 37501
rect 28533 37496 28580 37500
rect 28644 37498 28650 37500
rect 28901 37498 28967 37501
rect 31886 37498 31892 37500
rect 28533 37440 28538 37496
rect 28533 37436 28580 37440
rect 28644 37438 28690 37498
rect 28901 37496 31892 37498
rect 28901 37440 28906 37496
rect 28962 37440 31892 37496
rect 28901 37438 31892 37440
rect 28644 37436 28650 37438
rect 28533 37435 28599 37436
rect 28901 37435 28967 37438
rect 31886 37436 31892 37438
rect 31956 37436 31962 37500
rect 32305 37498 32371 37501
rect 32990 37498 32996 37500
rect 32305 37496 32996 37498
rect 32305 37440 32310 37496
rect 32366 37440 32996 37496
rect 32305 37438 32996 37440
rect 32305 37435 32371 37438
rect 32990 37436 32996 37438
rect 33060 37436 33066 37500
rect 33133 37498 33199 37501
rect 35433 37498 35499 37501
rect 33133 37496 35499 37498
rect 33133 37440 33138 37496
rect 33194 37440 35438 37496
rect 35494 37440 35499 37496
rect 33133 37438 35499 37440
rect 33133 37435 33199 37438
rect 35433 37435 35499 37438
rect 24710 37300 24716 37364
rect 24780 37362 24786 37364
rect 27838 37362 27844 37364
rect 24780 37302 27844 37362
rect 24780 37300 24786 37302
rect 27838 37300 27844 37302
rect 27908 37300 27914 37364
rect 28993 37362 29059 37365
rect 45870 37362 45876 37364
rect 28030 37302 28826 37362
rect 14406 37164 14412 37228
rect 14476 37226 14482 37228
rect 21081 37226 21147 37229
rect 14476 37224 21147 37226
rect 14476 37168 21086 37224
rect 21142 37168 21147 37224
rect 14476 37166 21147 37168
rect 14476 37164 14482 37166
rect 21081 37163 21147 37166
rect 22686 37164 22692 37228
rect 22756 37226 22762 37228
rect 23473 37226 23539 37229
rect 22756 37224 23539 37226
rect 22756 37168 23478 37224
rect 23534 37168 23539 37224
rect 22756 37166 23539 37168
rect 22756 37164 22762 37166
rect 23473 37163 23539 37166
rect 24894 37164 24900 37228
rect 24964 37226 24970 37228
rect 28030 37226 28090 37302
rect 24964 37166 28090 37226
rect 24964 37164 24970 37166
rect 28206 37164 28212 37228
rect 28276 37226 28282 37228
rect 28625 37226 28691 37229
rect 28276 37224 28691 37226
rect 28276 37168 28630 37224
rect 28686 37168 28691 37224
rect 28276 37166 28691 37168
rect 28766 37226 28826 37302
rect 28993 37360 45876 37362
rect 28993 37304 28998 37360
rect 29054 37304 45876 37360
rect 28993 37302 45876 37304
rect 28993 37299 29059 37302
rect 45870 37300 45876 37302
rect 45940 37300 45946 37364
rect 48405 37362 48471 37365
rect 53833 37362 53899 37365
rect 48405 37360 53899 37362
rect 48405 37304 48410 37360
rect 48466 37304 53838 37360
rect 53894 37304 53899 37360
rect 48405 37302 53899 37304
rect 48405 37299 48471 37302
rect 53833 37299 53899 37302
rect 37181 37226 37247 37229
rect 28766 37224 37247 37226
rect 28766 37168 37186 37224
rect 37242 37168 37247 37224
rect 28766 37166 37247 37168
rect 28276 37164 28282 37166
rect 28625 37163 28691 37166
rect 37181 37163 37247 37166
rect 12014 37028 12020 37092
rect 12084 37090 12090 37092
rect 21173 37090 21239 37093
rect 12084 37088 21239 37090
rect 12084 37032 21178 37088
rect 21234 37032 21239 37088
rect 12084 37030 21239 37032
rect 12084 37028 12090 37030
rect 21173 37027 21239 37030
rect 23606 37028 23612 37092
rect 23676 37090 23682 37092
rect 39389 37090 39455 37093
rect 23676 37088 39455 37090
rect 23676 37032 39394 37088
rect 39450 37032 39455 37088
rect 23676 37030 39455 37032
rect 23676 37028 23682 37030
rect 39389 37027 39455 37030
rect 1994 37024 2310 37025
rect 1994 36960 2000 37024
rect 2064 36960 2080 37024
rect 2144 36960 2160 37024
rect 2224 36960 2240 37024
rect 2304 36960 2310 37024
rect 1994 36959 2310 36960
rect 49994 37024 50310 37025
rect 49994 36960 50000 37024
rect 50064 36960 50080 37024
rect 50144 36960 50160 37024
rect 50224 36960 50240 37024
rect 50304 36960 50310 37024
rect 49994 36959 50310 36960
rect 64334 37024 64650 37025
rect 64334 36960 64340 37024
rect 64404 36960 64420 37024
rect 64484 36960 64500 37024
rect 64564 36960 64580 37024
rect 64644 36960 64650 37024
rect 64334 36959 64650 36960
rect 10910 36892 10916 36956
rect 10980 36954 10986 36956
rect 16205 36954 16271 36957
rect 10980 36952 16271 36954
rect 10980 36896 16210 36952
rect 16266 36896 16271 36952
rect 10980 36894 16271 36896
rect 10980 36892 10986 36894
rect 16205 36891 16271 36894
rect 19333 36954 19399 36957
rect 38878 36954 38884 36956
rect 19333 36952 38884 36954
rect 19333 36896 19338 36952
rect 19394 36896 38884 36952
rect 19333 36894 38884 36896
rect 19333 36891 19399 36894
rect 38878 36892 38884 36894
rect 38948 36892 38954 36956
rect 9622 36756 9628 36820
rect 9692 36818 9698 36820
rect 20713 36818 20779 36821
rect 9692 36816 20779 36818
rect 9692 36760 20718 36816
rect 20774 36760 20779 36816
rect 9692 36758 20779 36760
rect 9692 36756 9698 36758
rect 20713 36755 20779 36758
rect 23197 36818 23263 36821
rect 37590 36818 37596 36820
rect 23197 36816 37596 36818
rect 23197 36760 23202 36816
rect 23258 36760 37596 36816
rect 23197 36758 37596 36760
rect 23197 36755 23263 36758
rect 37590 36756 37596 36758
rect 37660 36756 37666 36820
rect 37733 36818 37799 36821
rect 62614 36818 62620 36820
rect 37733 36816 62620 36818
rect 37733 36760 37738 36816
rect 37794 36760 62620 36816
rect 37733 36758 62620 36760
rect 37733 36755 37799 36758
rect 62614 36756 62620 36758
rect 62684 36756 62690 36820
rect 5022 36620 5028 36684
rect 5092 36682 5098 36684
rect 12341 36682 12407 36685
rect 5092 36680 12407 36682
rect 5092 36624 12346 36680
rect 12402 36624 12407 36680
rect 5092 36622 12407 36624
rect 5092 36620 5098 36622
rect 12341 36619 12407 36622
rect 16389 36682 16455 36685
rect 39982 36682 39988 36684
rect 16389 36680 39988 36682
rect 16389 36624 16394 36680
rect 16450 36624 39988 36680
rect 16389 36622 39988 36624
rect 16389 36619 16455 36622
rect 39982 36620 39988 36622
rect 40052 36620 40058 36684
rect 41689 36682 41755 36685
rect 65609 36682 65675 36685
rect 41689 36680 65675 36682
rect 41689 36624 41694 36680
rect 41750 36624 65614 36680
rect 65670 36624 65675 36680
rect 41689 36622 65675 36624
rect 41689 36619 41755 36622
rect 65609 36619 65675 36622
rect 6126 36484 6132 36548
rect 6196 36546 6202 36548
rect 17953 36546 18019 36549
rect 6196 36544 18019 36546
rect 6196 36488 17958 36544
rect 18014 36488 18019 36544
rect 6196 36486 18019 36488
rect 6196 36484 6202 36486
rect 17953 36483 18019 36486
rect 26734 36484 26740 36548
rect 26804 36546 26810 36548
rect 27521 36546 27587 36549
rect 26804 36544 27587 36546
rect 26804 36488 27526 36544
rect 27582 36488 27587 36544
rect 26804 36486 27587 36488
rect 26804 36484 26810 36486
rect 27521 36483 27587 36486
rect 36537 36546 36603 36549
rect 63309 36546 63375 36549
rect 36537 36544 63375 36546
rect 36537 36488 36542 36544
rect 36598 36488 63314 36544
rect 63370 36488 63375 36544
rect 36537 36486 63375 36488
rect 36537 36483 36603 36486
rect 63309 36483 63375 36486
rect 65254 36480 65570 36481
rect 65254 36416 65260 36480
rect 65324 36416 65340 36480
rect 65404 36416 65420 36480
rect 65484 36416 65500 36480
rect 65564 36416 65570 36480
rect 65254 36415 65570 36416
rect 22502 36348 22508 36412
rect 22572 36410 22578 36412
rect 27245 36410 27311 36413
rect 22572 36408 27311 36410
rect 22572 36352 27250 36408
rect 27306 36352 27311 36408
rect 22572 36350 27311 36352
rect 22572 36348 22578 36350
rect 27245 36347 27311 36350
rect 33174 36348 33180 36412
rect 33244 36410 33250 36412
rect 42701 36410 42767 36413
rect 33244 36408 42767 36410
rect 33244 36352 42706 36408
rect 42762 36352 42767 36408
rect 33244 36350 42767 36352
rect 33244 36348 33250 36350
rect 42701 36347 42767 36350
rect 21582 36212 21588 36276
rect 21652 36274 21658 36276
rect 27613 36274 27679 36277
rect 35525 36274 35591 36277
rect 21652 36272 27679 36274
rect 21652 36216 27618 36272
rect 27674 36216 27679 36272
rect 21652 36214 27679 36216
rect 21652 36212 21658 36214
rect 27613 36211 27679 36214
rect 27846 36272 35591 36274
rect 27846 36216 35530 36272
rect 35586 36216 35591 36272
rect 27846 36214 35591 36216
rect 16614 36076 16620 36140
rect 16684 36138 16690 36140
rect 25405 36138 25471 36141
rect 16684 36136 25471 36138
rect 16684 36080 25410 36136
rect 25466 36080 25471 36136
rect 16684 36078 25471 36080
rect 16684 36076 16690 36078
rect 25405 36075 25471 36078
rect 13152 35940 13158 36004
rect 13222 36002 13228 36004
rect 17861 36002 17927 36005
rect 20989 36002 21055 36005
rect 24669 36004 24735 36005
rect 13222 36000 17927 36002
rect 13222 35944 17866 36000
rect 17922 35944 17927 36000
rect 13222 35942 17927 35944
rect 13222 35940 13228 35942
rect 17861 35939 17927 35942
rect 19198 36000 21055 36002
rect 19198 35944 20994 36000
rect 21050 35944 21055 36000
rect 19198 35942 21055 35944
rect 17824 35804 17830 35868
rect 17894 35866 17900 35868
rect 19198 35866 19258 35942
rect 20989 35939 21055 35942
rect 22970 35942 23490 36002
rect 17894 35806 19258 35866
rect 17894 35804 17900 35806
rect 19466 35804 19472 35868
rect 19536 35866 19542 35868
rect 20621 35866 20687 35869
rect 19536 35864 20687 35866
rect 19536 35808 20626 35864
rect 20682 35808 20687 35864
rect 19536 35806 20687 35808
rect 19536 35804 19542 35806
rect 20621 35803 20687 35806
rect 20962 35804 20968 35868
rect 21032 35866 21038 35868
rect 22970 35866 23030 35942
rect 23197 35868 23263 35869
rect 23192 35866 23198 35868
rect 21032 35806 23030 35866
rect 23110 35806 23198 35866
rect 21032 35804 21038 35806
rect 23192 35804 23198 35806
rect 23262 35804 23268 35868
rect 23430 35866 23490 35942
rect 24669 36000 24692 36004
rect 24756 36002 24762 36004
rect 24669 35944 24674 36000
rect 24669 35940 24692 35944
rect 24756 35942 24826 36002
rect 24756 35940 24762 35942
rect 26458 35940 26464 36004
rect 26528 36002 26534 36004
rect 27846 36002 27906 36214
rect 35525 36211 35591 36214
rect 38653 36274 38719 36277
rect 62757 36274 62823 36277
rect 38653 36272 62823 36274
rect 38653 36216 38658 36272
rect 38714 36216 62762 36272
rect 62818 36216 62823 36272
rect 38653 36214 62823 36216
rect 38653 36211 38719 36214
rect 62757 36211 62823 36214
rect 33409 36138 33475 36141
rect 29200 36136 33475 36138
rect 29200 36080 33414 36136
rect 33470 36080 33475 36136
rect 29200 36078 33475 36080
rect 29200 36004 29260 36078
rect 33409 36075 33475 36078
rect 38653 36138 38719 36141
rect 63493 36138 63559 36141
rect 38653 36136 63559 36138
rect 38653 36080 38658 36136
rect 38714 36080 63498 36136
rect 63554 36080 63559 36136
rect 38653 36078 63559 36080
rect 38653 36075 38719 36078
rect 63493 36075 63559 36078
rect 30649 36004 30715 36005
rect 26528 35942 27906 36002
rect 26528 35940 26534 35942
rect 29192 35940 29198 36004
rect 29262 35940 29268 36004
rect 30649 36002 30678 36004
rect 30054 35942 30482 36002
rect 30586 36000 30678 36002
rect 30586 35944 30654 36000
rect 30586 35942 30678 35944
rect 24669 35939 24735 35940
rect 25497 35866 25563 35869
rect 25865 35868 25931 35869
rect 23430 35864 25563 35866
rect 23430 35808 25502 35864
rect 25558 35808 25563 35864
rect 23430 35806 25563 35808
rect 23197 35803 23263 35804
rect 25497 35803 25563 35806
rect 25862 35804 25868 35868
rect 25932 35866 25938 35868
rect 25932 35806 26022 35866
rect 25932 35804 25938 35806
rect 29504 35804 29510 35868
rect 29574 35866 29580 35868
rect 30054 35866 30114 35942
rect 30281 35868 30347 35869
rect 30230 35866 30236 35868
rect 29574 35806 30114 35866
rect 30190 35806 30236 35866
rect 30300 35864 30347 35868
rect 30342 35808 30347 35864
rect 29574 35804 29580 35806
rect 30230 35804 30236 35806
rect 30300 35804 30347 35808
rect 30422 35866 30482 35942
rect 30649 35940 30678 35942
rect 30742 35940 30748 36004
rect 30925 36002 30991 36005
rect 31192 36002 31198 36004
rect 30925 36000 31198 36002
rect 30925 35944 30930 36000
rect 30986 35944 31198 36000
rect 30925 35942 31198 35944
rect 30649 35939 30715 35940
rect 30925 35939 30991 35942
rect 31192 35940 31198 35942
rect 31262 35940 31268 36004
rect 31702 35940 31708 36004
rect 31772 36002 31778 36004
rect 32070 36002 32076 36004
rect 31772 35942 32076 36002
rect 31772 35940 31778 35942
rect 32070 35940 32076 35942
rect 32140 35940 32146 36004
rect 35801 36002 35867 36005
rect 63769 36002 63835 36005
rect 64086 36002 64092 36004
rect 35801 36000 62130 36002
rect 35801 35944 35806 36000
rect 35862 35944 62130 36000
rect 35801 35942 62130 35944
rect 35801 35939 35867 35942
rect 31661 35866 31727 35869
rect 30422 35864 31727 35866
rect 30422 35808 31666 35864
rect 31722 35808 31727 35864
rect 30422 35806 31727 35808
rect 25865 35803 25931 35804
rect 30281 35803 30347 35804
rect 31661 35803 31727 35806
rect 33910 35804 33916 35868
rect 33980 35866 33986 35868
rect 34145 35866 34211 35869
rect 33980 35864 34211 35866
rect 33980 35808 34150 35864
rect 34206 35808 34211 35864
rect 33980 35806 34211 35808
rect 33980 35804 33986 35806
rect 34145 35803 34211 35806
rect 34421 35866 34487 35869
rect 36512 35866 36518 35868
rect 34421 35864 36518 35866
rect 34421 35808 34426 35864
rect 34482 35808 36518 35864
rect 34421 35806 36518 35808
rect 34421 35803 34487 35806
rect 36512 35804 36518 35806
rect 36582 35804 36588 35868
rect 40125 35866 40191 35869
rect 43529 35868 43595 35869
rect 42352 35866 42358 35868
rect 40125 35864 42358 35866
rect 40125 35808 40130 35864
rect 40186 35808 42358 35864
rect 40125 35806 42358 35808
rect 40125 35803 40191 35806
rect 42352 35804 42358 35806
rect 42422 35804 42428 35868
rect 43520 35866 43526 35868
rect 43438 35806 43526 35866
rect 43520 35804 43526 35806
rect 43590 35804 43596 35868
rect 62070 35866 62130 35942
rect 63769 36000 64092 36002
rect 63769 35944 63774 36000
rect 63830 35944 64092 36000
rect 63769 35942 64092 35944
rect 63769 35939 63835 35942
rect 64086 35940 64092 35942
rect 64156 35940 64162 36004
rect 64334 35936 64650 35937
rect 64334 35872 64340 35936
rect 64404 35872 64420 35936
rect 64484 35872 64500 35936
rect 64564 35872 64580 35936
rect 64644 35872 64650 35936
rect 64334 35871 64650 35872
rect 63534 35866 63540 35868
rect 62070 35806 63540 35866
rect 63534 35804 63540 35806
rect 63604 35804 63610 35868
rect 43529 35803 43595 35804
rect 7322 35668 7328 35732
rect 7392 35730 7398 35732
rect 8201 35730 8267 35733
rect 7392 35728 8267 35730
rect 7392 35672 8206 35728
rect 8262 35672 8267 35728
rect 7392 35670 8267 35672
rect 7392 35668 7398 35670
rect 8201 35667 8267 35670
rect 8477 35732 8543 35733
rect 20069 35732 20135 35733
rect 8477 35728 8486 35732
rect 8550 35730 8556 35732
rect 20022 35730 20028 35732
rect 8477 35672 8482 35728
rect 8477 35668 8486 35672
rect 8550 35670 8634 35730
rect 19978 35670 20028 35730
rect 20092 35728 20135 35732
rect 20130 35672 20135 35728
rect 8550 35668 8556 35670
rect 20022 35668 20028 35670
rect 20092 35668 20135 35672
rect 8477 35667 8543 35668
rect 20069 35667 20135 35668
rect 21173 35732 21239 35733
rect 22001 35732 22067 35733
rect 22185 35732 22251 35733
rect 23013 35732 23079 35733
rect 23565 35732 23631 35733
rect 30005 35732 30071 35733
rect 21173 35728 21196 35732
rect 21260 35730 21266 35732
rect 21962 35730 21968 35732
rect 21173 35672 21178 35728
rect 21173 35668 21196 35672
rect 21260 35670 21330 35730
rect 21910 35670 21968 35730
rect 22032 35728 22067 35732
rect 22062 35672 22067 35728
rect 21260 35668 21266 35670
rect 21962 35668 21968 35670
rect 22032 35668 22067 35672
rect 22134 35668 22140 35732
rect 22204 35730 22251 35732
rect 22962 35730 22968 35732
rect 22204 35728 22296 35730
rect 22246 35672 22296 35728
rect 22204 35670 22296 35672
rect 22922 35670 22968 35730
rect 23032 35728 23079 35732
rect 23526 35730 23532 35732
rect 23074 35672 23079 35728
rect 22204 35668 22251 35670
rect 22962 35668 22968 35670
rect 23032 35668 23079 35672
rect 23474 35670 23532 35730
rect 23596 35728 23631 35732
rect 23626 35672 23631 35728
rect 23526 35668 23532 35670
rect 23596 35668 23631 35672
rect 25204 35668 25210 35732
rect 25274 35730 25280 35732
rect 26182 35730 26188 35732
rect 25274 35670 26188 35730
rect 25274 35668 25280 35670
rect 26182 35668 26188 35670
rect 26252 35668 26258 35732
rect 29962 35730 29968 35732
rect 29914 35670 29968 35730
rect 30032 35728 30071 35732
rect 30066 35672 30071 35728
rect 29962 35668 29968 35670
rect 30032 35668 30071 35672
rect 21173 35667 21239 35668
rect 22001 35667 22067 35668
rect 22185 35667 22251 35668
rect 23013 35667 23079 35668
rect 23565 35667 23631 35668
rect 30005 35667 30071 35668
rect 31017 35730 31083 35733
rect 32870 35730 32876 35732
rect 31017 35728 32876 35730
rect 31017 35672 31022 35728
rect 31078 35672 32876 35728
rect 31017 35670 32876 35672
rect 31017 35667 31083 35670
rect 32870 35668 32876 35670
rect 32940 35668 32946 35732
rect 33133 35730 33199 35733
rect 33450 35730 33456 35732
rect 33133 35728 33456 35730
rect 33133 35672 33138 35728
rect 33194 35672 33456 35728
rect 33133 35670 33456 35672
rect 33133 35667 33199 35670
rect 33450 35668 33456 35670
rect 33520 35668 33526 35732
rect 33593 35730 33659 35733
rect 33726 35730 33732 35732
rect 33593 35728 33732 35730
rect 33593 35672 33598 35728
rect 33654 35672 33732 35728
rect 33593 35670 33732 35672
rect 33593 35667 33659 35670
rect 33726 35668 33732 35670
rect 33796 35668 33802 35732
rect 40033 35730 40099 35733
rect 41178 35730 41184 35732
rect 40033 35728 41184 35730
rect 40033 35672 40038 35728
rect 40094 35672 41184 35728
rect 40033 35670 41184 35672
rect 40033 35667 40099 35670
rect 41178 35668 41184 35670
rect 41248 35668 41254 35732
rect 42701 35730 42767 35733
rect 44674 35730 44680 35732
rect 42701 35728 44680 35730
rect 42701 35672 42706 35728
rect 42762 35672 44680 35728
rect 42701 35670 44680 35672
rect 42701 35667 42767 35670
rect 44674 35668 44680 35670
rect 44744 35668 44750 35732
rect 56041 35730 56107 35733
rect 56240 35730 56246 35732
rect 56041 35728 56246 35730
rect 56041 35672 56046 35728
rect 56102 35672 56246 35728
rect 56041 35670 56246 35672
rect 56041 35667 56107 35670
rect 56240 35668 56246 35670
rect 56310 35730 56316 35732
rect 63861 35730 63927 35733
rect 56310 35728 63927 35730
rect 56310 35672 63866 35728
rect 63922 35672 63927 35728
rect 56310 35670 63927 35672
rect 56310 35668 56316 35670
rect 63861 35667 63927 35670
rect 62798 35532 62804 35596
rect 62868 35594 62874 35596
rect 63585 35594 63651 35597
rect 62868 35592 63651 35594
rect 62868 35536 63590 35592
rect 63646 35536 63651 35592
rect 62868 35534 63651 35536
rect 62868 35532 62874 35534
rect 63585 35531 63651 35534
rect 400 35492 748 35514
rect 400 35428 422 35492
rect 486 35428 502 35492
rect 566 35428 582 35492
rect 646 35428 662 35492
rect 726 35428 748 35492
rect 400 35412 748 35428
rect 400 35348 422 35412
rect 486 35348 502 35412
rect 566 35348 582 35412
rect 646 35348 662 35412
rect 726 35348 748 35412
rect 400 35332 748 35348
rect 400 35268 422 35332
rect 486 35268 502 35332
rect 566 35268 582 35332
rect 646 35268 662 35332
rect 726 35268 748 35332
rect 400 35252 748 35268
rect 400 35188 422 35252
rect 486 35188 502 35252
rect 566 35188 582 35252
rect 646 35188 662 35252
rect 726 35188 748 35252
rect 400 35166 748 35188
rect 1992 35492 2312 35514
rect 1992 35428 2000 35492
rect 2064 35428 2080 35492
rect 2144 35428 2160 35492
rect 2224 35428 2240 35492
rect 2304 35428 2312 35492
rect 1992 35412 2312 35428
rect 1992 35348 2000 35412
rect 2064 35348 2080 35412
rect 2144 35348 2160 35412
rect 2224 35348 2240 35412
rect 2304 35348 2312 35412
rect 1992 35332 2312 35348
rect 1992 35268 2000 35332
rect 2064 35268 2080 35332
rect 2144 35268 2160 35332
rect 2224 35268 2240 35332
rect 2304 35268 2312 35332
rect 1992 35252 2312 35268
rect 1992 35188 2000 35252
rect 2064 35188 2080 35252
rect 2144 35188 2160 35252
rect 2224 35188 2240 35252
rect 2304 35188 2312 35252
rect 1992 35166 2312 35188
rect 49992 35492 50312 35514
rect 49992 35428 50000 35492
rect 50064 35428 50080 35492
rect 50144 35428 50160 35492
rect 50224 35428 50240 35492
rect 50304 35428 50312 35492
rect 49992 35412 50312 35428
rect 49992 35348 50000 35412
rect 50064 35348 50080 35412
rect 50144 35348 50160 35412
rect 50224 35348 50240 35412
rect 50304 35348 50312 35412
rect 49992 35332 50312 35348
rect 49992 35268 50000 35332
rect 50064 35268 50080 35332
rect 50144 35268 50160 35332
rect 50224 35268 50240 35332
rect 50304 35268 50312 35332
rect 49992 35252 50312 35268
rect 49992 35188 50000 35252
rect 50064 35188 50080 35252
rect 50144 35188 50160 35252
rect 50224 35188 50240 35252
rect 50304 35188 50312 35252
rect 49992 35166 50312 35188
rect 62188 35492 62536 35514
rect 62188 35428 62210 35492
rect 62274 35428 62290 35492
rect 62354 35428 62370 35492
rect 62434 35428 62450 35492
rect 62514 35428 62536 35492
rect 62188 35412 62536 35428
rect 62188 35348 62210 35412
rect 62274 35348 62290 35412
rect 62354 35348 62370 35412
rect 62434 35348 62450 35412
rect 62514 35348 62536 35412
rect 62188 35332 62536 35348
rect 62188 35268 62210 35332
rect 62274 35268 62290 35332
rect 62354 35268 62370 35332
rect 62434 35268 62450 35332
rect 62514 35268 62536 35332
rect 65254 35392 65570 35393
rect 65254 35328 65260 35392
rect 65324 35328 65340 35392
rect 65404 35328 65420 35392
rect 65484 35328 65500 35392
rect 65564 35328 65570 35392
rect 65254 35327 65570 35328
rect 62188 35252 62536 35268
rect 62188 35188 62210 35252
rect 62274 35188 62290 35252
rect 62354 35188 62370 35252
rect 62434 35188 62450 35252
rect 62514 35188 62536 35252
rect 62188 35166 62536 35188
rect 62573 35050 62639 35053
rect 63718 35050 63724 35052
rect 62573 35048 63724 35050
rect 62573 34992 62578 35048
rect 62634 34992 63724 35048
rect 62573 34990 63724 34992
rect 62573 34987 62639 34990
rect 63718 34988 63724 34990
rect 63788 34988 63794 35052
rect 64334 34848 64650 34849
rect 1096 34796 1444 34818
rect 1096 34732 1118 34796
rect 1182 34732 1198 34796
rect 1262 34732 1278 34796
rect 1342 34732 1358 34796
rect 1422 34732 1444 34796
rect 1096 34716 1444 34732
rect 1096 34652 1118 34716
rect 1182 34652 1198 34716
rect 1262 34652 1278 34716
rect 1342 34652 1358 34716
rect 1422 34652 1444 34716
rect 1096 34636 1444 34652
rect 1096 34572 1118 34636
rect 1182 34572 1198 34636
rect 1262 34572 1278 34636
rect 1342 34572 1358 34636
rect 1422 34572 1444 34636
rect 1096 34556 1444 34572
rect 1096 34492 1118 34556
rect 1182 34492 1198 34556
rect 1262 34492 1278 34556
rect 1342 34492 1358 34556
rect 1422 34492 1444 34556
rect 1096 34470 1444 34492
rect 2912 34796 3232 34818
rect 2912 34732 2920 34796
rect 2984 34732 3000 34796
rect 3064 34732 3080 34796
rect 3144 34732 3160 34796
rect 3224 34732 3232 34796
rect 2912 34716 3232 34732
rect 2912 34652 2920 34716
rect 2984 34652 3000 34716
rect 3064 34652 3080 34716
rect 3144 34652 3160 34716
rect 3224 34652 3232 34716
rect 2912 34636 3232 34652
rect 2912 34572 2920 34636
rect 2984 34572 3000 34636
rect 3064 34572 3080 34636
rect 3144 34572 3160 34636
rect 3224 34572 3232 34636
rect 2912 34556 3232 34572
rect 2912 34492 2920 34556
rect 2984 34492 3000 34556
rect 3064 34492 3080 34556
rect 3144 34492 3160 34556
rect 3224 34492 3232 34556
rect 2912 34470 3232 34492
rect 50912 34796 51232 34818
rect 50912 34732 50920 34796
rect 50984 34732 51000 34796
rect 51064 34732 51080 34796
rect 51144 34732 51160 34796
rect 51224 34732 51232 34796
rect 50912 34716 51232 34732
rect 50912 34652 50920 34716
rect 50984 34652 51000 34716
rect 51064 34652 51080 34716
rect 51144 34652 51160 34716
rect 51224 34652 51232 34716
rect 50912 34636 51232 34652
rect 50912 34572 50920 34636
rect 50984 34572 51000 34636
rect 51064 34572 51080 34636
rect 51144 34572 51160 34636
rect 51224 34572 51232 34636
rect 50912 34556 51232 34572
rect 50912 34492 50920 34556
rect 50984 34492 51000 34556
rect 51064 34492 51080 34556
rect 51144 34492 51160 34556
rect 51224 34492 51232 34556
rect 50912 34470 51232 34492
rect 61492 34796 61840 34818
rect 61492 34732 61514 34796
rect 61578 34732 61594 34796
rect 61658 34732 61674 34796
rect 61738 34732 61754 34796
rect 61818 34732 61840 34796
rect 64334 34784 64340 34848
rect 64404 34784 64420 34848
rect 64484 34784 64500 34848
rect 64564 34784 64580 34848
rect 64644 34784 64650 34848
rect 64334 34783 64650 34784
rect 61492 34716 61840 34732
rect 61492 34652 61514 34716
rect 61578 34652 61594 34716
rect 61658 34652 61674 34716
rect 61738 34652 61754 34716
rect 61818 34652 61840 34716
rect 61492 34636 61840 34652
rect 61492 34572 61514 34636
rect 61578 34572 61594 34636
rect 61658 34572 61674 34636
rect 61738 34572 61754 34636
rect 61818 34572 61840 34636
rect 61492 34556 61840 34572
rect 61492 34492 61514 34556
rect 61578 34492 61594 34556
rect 61658 34492 61674 34556
rect 61738 34492 61754 34556
rect 61818 34492 61840 34556
rect 61492 34470 61840 34492
rect 65254 34304 65570 34305
rect 65254 34240 65260 34304
rect 65324 34240 65340 34304
rect 65404 34240 65420 34304
rect 65484 34240 65500 34304
rect 65564 34240 65570 34304
rect 65254 34239 65570 34240
rect 64334 33760 64650 33761
rect 64334 33696 64340 33760
rect 64404 33696 64420 33760
rect 64484 33696 64500 33760
rect 64564 33696 64580 33760
rect 64644 33696 64650 33760
rect 64334 33695 64650 33696
rect 65254 33216 65570 33217
rect 65254 33152 65260 33216
rect 65324 33152 65340 33216
rect 65404 33152 65420 33216
rect 65484 33152 65500 33216
rect 65564 33152 65570 33216
rect 65254 33151 65570 33152
rect 63493 33146 63559 33149
rect 63902 33146 63908 33148
rect 63493 33144 63908 33146
rect 63493 33088 63498 33144
rect 63554 33088 63908 33144
rect 63493 33086 63908 33088
rect 63493 33083 63559 33086
rect 63902 33084 63908 33086
rect 63972 33084 63978 33148
rect 64334 32672 64650 32673
rect 64334 32608 64340 32672
rect 64404 32608 64420 32672
rect 64484 32608 64500 32672
rect 64564 32608 64580 32672
rect 64644 32608 64650 32672
rect 64334 32607 64650 32608
rect 64086 32404 64092 32468
rect 64156 32466 64162 32468
rect 64689 32466 64755 32469
rect 64156 32464 64755 32466
rect 64156 32408 64694 32464
rect 64750 32408 64755 32464
rect 64156 32406 64755 32408
rect 64156 32404 64162 32406
rect 64689 32403 64755 32406
rect 65254 32128 65570 32129
rect 65254 32064 65260 32128
rect 65324 32064 65340 32128
rect 65404 32064 65420 32128
rect 65484 32064 65500 32128
rect 65564 32064 65570 32128
rect 65254 32063 65570 32064
rect 66161 31920 66227 31925
rect 66161 31864 66166 31920
rect 66222 31864 66227 31920
rect 66161 31859 66227 31864
rect 64965 31786 65031 31789
rect 65333 31786 65399 31789
rect 64965 31784 65399 31786
rect 64965 31728 64970 31784
rect 65026 31728 65338 31784
rect 65394 31728 65399 31784
rect 64965 31726 65399 31728
rect 64965 31723 65031 31726
rect 65333 31723 65399 31726
rect 65885 31786 65951 31789
rect 66164 31786 66224 31859
rect 65885 31784 66224 31786
rect 65885 31728 65890 31784
rect 65946 31728 66224 31784
rect 65885 31726 66224 31728
rect 65885 31723 65951 31726
rect 64334 31584 64650 31585
rect 64334 31520 64340 31584
rect 64404 31520 64420 31584
rect 64484 31520 64500 31584
rect 64564 31520 64580 31584
rect 64644 31520 64650 31584
rect 64334 31519 64650 31520
rect 65254 31040 65570 31041
rect 65254 30976 65260 31040
rect 65324 30976 65340 31040
rect 65404 30976 65420 31040
rect 65484 30976 65500 31040
rect 65564 30976 65570 31040
rect 65254 30975 65570 30976
rect 62665 30940 62731 30943
rect 62504 30938 62731 30940
rect 62504 30882 62670 30938
rect 62726 30882 62731 30938
rect 62504 30880 62731 30882
rect 62665 30877 62731 30880
rect 64334 30496 64650 30497
rect 64334 30432 64340 30496
rect 64404 30432 64420 30496
rect 64484 30432 64500 30496
rect 64564 30432 64580 30496
rect 64644 30432 64650 30496
rect 64334 30431 64650 30432
rect 65254 29952 65570 29953
rect 65254 29888 65260 29952
rect 65324 29888 65340 29952
rect 65404 29888 65420 29952
rect 65484 29888 65500 29952
rect 65564 29888 65570 29952
rect 65254 29887 65570 29888
rect 64334 29408 64650 29409
rect 64334 29344 64340 29408
rect 64404 29344 64420 29408
rect 64484 29344 64500 29408
rect 64564 29344 64580 29408
rect 64644 29344 64650 29408
rect 64334 29343 64650 29344
rect 62757 29240 62823 29243
rect 62504 29238 62823 29240
rect 62504 29182 62762 29238
rect 62818 29182 62823 29238
rect 62504 29180 62823 29182
rect 62757 29177 62823 29180
rect 65254 28864 65570 28865
rect 65254 28800 65260 28864
rect 65324 28800 65340 28864
rect 65404 28800 65420 28864
rect 65484 28800 65500 28864
rect 65564 28800 65570 28864
rect 65254 28799 65570 28800
rect 64334 28320 64650 28321
rect 64334 28256 64340 28320
rect 64404 28256 64420 28320
rect 64484 28256 64500 28320
rect 64564 28256 64580 28320
rect 64644 28256 64650 28320
rect 64334 28255 64650 28256
rect 65254 27776 65570 27777
rect 65254 27712 65260 27776
rect 65324 27712 65340 27776
rect 65404 27712 65420 27776
rect 65484 27712 65500 27776
rect 65564 27712 65570 27776
rect 65254 27711 65570 27712
rect 64334 27232 64650 27233
rect 64334 27168 64340 27232
rect 64404 27168 64420 27232
rect 64484 27168 64500 27232
rect 64564 27168 64580 27232
rect 64644 27168 64650 27232
rect 64334 27167 64650 27168
rect 65254 26688 65570 26689
rect 65254 26624 65260 26688
rect 65324 26624 65340 26688
rect 65404 26624 65420 26688
rect 65484 26624 65500 26688
rect 65564 26624 65570 26688
rect 65254 26623 65570 26624
rect 64334 26144 64650 26145
rect 64334 26080 64340 26144
rect 64404 26080 64420 26144
rect 64484 26080 64500 26144
rect 64564 26080 64580 26144
rect 64644 26080 64650 26144
rect 64334 26079 64650 26080
rect 65254 25600 65570 25601
rect 65254 25536 65260 25600
rect 65324 25536 65340 25600
rect 65404 25536 65420 25600
rect 65484 25536 65500 25600
rect 65564 25536 65570 25600
rect 65254 25535 65570 25536
rect 64334 25056 64650 25057
rect 64334 24992 64340 25056
rect 64404 24992 64420 25056
rect 64484 24992 64500 25056
rect 64564 24992 64580 25056
rect 64644 24992 64650 25056
rect 64334 24991 64650 24992
rect 65254 24512 65570 24513
rect 65254 24448 65260 24512
rect 65324 24448 65340 24512
rect 65404 24448 65420 24512
rect 65484 24448 65500 24512
rect 65564 24448 65570 24512
rect 65254 24447 65570 24448
rect 64334 23968 64650 23969
rect 64334 23904 64340 23968
rect 64404 23904 64420 23968
rect 64484 23904 64500 23968
rect 64564 23904 64580 23968
rect 64644 23904 64650 23968
rect 64334 23903 64650 23904
rect 65254 23424 65570 23425
rect 65254 23360 65260 23424
rect 65324 23360 65340 23424
rect 65404 23360 65420 23424
rect 65484 23360 65500 23424
rect 65564 23360 65570 23424
rect 65254 23359 65570 23360
rect 64334 22880 64650 22881
rect 64334 22816 64340 22880
rect 64404 22816 64420 22880
rect 64484 22816 64500 22880
rect 64564 22816 64580 22880
rect 64644 22816 64650 22880
rect 64334 22815 64650 22816
rect 65254 22336 65570 22337
rect 65254 22272 65260 22336
rect 65324 22272 65340 22336
rect 65404 22272 65420 22336
rect 65484 22272 65500 22336
rect 65564 22272 65570 22336
rect 65254 22271 65570 22272
rect 64334 21792 64650 21793
rect 64334 21728 64340 21792
rect 64404 21728 64420 21792
rect 64484 21728 64500 21792
rect 64564 21728 64580 21792
rect 64644 21728 64650 21792
rect 64334 21727 64650 21728
rect 65254 21248 65570 21249
rect 65254 21184 65260 21248
rect 65324 21184 65340 21248
rect 65404 21184 65420 21248
rect 65484 21184 65500 21248
rect 65564 21184 65570 21248
rect 65254 21183 65570 21184
rect 64334 20704 64650 20705
rect 64334 20640 64340 20704
rect 64404 20640 64420 20704
rect 64484 20640 64500 20704
rect 64564 20640 64580 20704
rect 64644 20640 64650 20704
rect 64334 20639 64650 20640
rect 65254 20160 65570 20161
rect 65254 20096 65260 20160
rect 65324 20096 65340 20160
rect 65404 20096 65420 20160
rect 65484 20096 65500 20160
rect 65564 20096 65570 20160
rect 65254 20095 65570 20096
rect 64334 19616 64650 19617
rect 64334 19552 64340 19616
rect 64404 19552 64420 19616
rect 64484 19552 64500 19616
rect 64564 19552 64580 19616
rect 64644 19552 64650 19616
rect 64334 19551 64650 19552
rect 65254 19072 65570 19073
rect 65254 19008 65260 19072
rect 65324 19008 65340 19072
rect 65404 19008 65420 19072
rect 65484 19008 65500 19072
rect 65564 19008 65570 19072
rect 65254 19007 65570 19008
rect 64334 18528 64650 18529
rect 64334 18464 64340 18528
rect 64404 18464 64420 18528
rect 64484 18464 64500 18528
rect 64564 18464 64580 18528
rect 64644 18464 64650 18528
rect 64334 18463 64650 18464
rect 65254 17984 65570 17985
rect 65254 17920 65260 17984
rect 65324 17920 65340 17984
rect 65404 17920 65420 17984
rect 65484 17920 65500 17984
rect 65564 17920 65570 17984
rect 65254 17919 65570 17920
rect 63718 17852 63724 17916
rect 63788 17914 63794 17916
rect 64689 17914 64755 17917
rect 63788 17912 64755 17914
rect 63788 17856 64694 17912
rect 64750 17856 64755 17912
rect 63788 17854 64755 17856
rect 63788 17852 63794 17854
rect 64689 17851 64755 17854
rect 64334 17440 64650 17441
rect 64334 17376 64340 17440
rect 64404 17376 64420 17440
rect 64484 17376 64500 17440
rect 64564 17376 64580 17440
rect 64644 17376 64650 17440
rect 64334 17375 64650 17376
rect 62573 17234 62639 17237
rect 62798 17234 62804 17236
rect 62573 17232 62804 17234
rect 62573 17176 62578 17232
rect 62634 17176 62804 17232
rect 62573 17174 62804 17176
rect 62573 17171 62639 17174
rect 62798 17172 62804 17174
rect 62868 17172 62874 17236
rect 65254 16896 65570 16897
rect 65254 16832 65260 16896
rect 65324 16832 65340 16896
rect 65404 16832 65420 16896
rect 65484 16832 65500 16896
rect 65564 16832 65570 16896
rect 65254 16831 65570 16832
rect 64334 16352 64650 16353
rect 64334 16288 64340 16352
rect 64404 16288 64420 16352
rect 64484 16288 64500 16352
rect 64564 16288 64580 16352
rect 64644 16288 64650 16352
rect 64334 16287 64650 16288
rect 65254 15808 65570 15809
rect 65254 15744 65260 15808
rect 65324 15744 65340 15808
rect 65404 15744 65420 15808
rect 65484 15744 65500 15808
rect 65564 15744 65570 15808
rect 65254 15743 65570 15744
rect 62614 15676 62620 15740
rect 62684 15738 62690 15740
rect 64781 15738 64847 15741
rect 62684 15736 64847 15738
rect 62684 15680 64786 15736
rect 64842 15680 64847 15736
rect 62684 15678 64847 15680
rect 62684 15676 62690 15678
rect 64781 15675 64847 15678
rect 64334 15264 64650 15265
rect 64334 15200 64340 15264
rect 64404 15200 64420 15264
rect 64484 15200 64500 15264
rect 64564 15200 64580 15264
rect 64644 15200 64650 15264
rect 64334 15199 64650 15200
rect 65254 14720 65570 14721
rect 65254 14656 65260 14720
rect 65324 14656 65340 14720
rect 65404 14656 65420 14720
rect 65484 14656 65500 14720
rect 65564 14656 65570 14720
rect 65254 14655 65570 14656
rect 64334 14176 64650 14177
rect 64334 14112 64340 14176
rect 64404 14112 64420 14176
rect 64484 14112 64500 14176
rect 64564 14112 64580 14176
rect 64644 14112 64650 14176
rect 64334 14111 64650 14112
rect 65254 13632 65570 13633
rect 65254 13568 65260 13632
rect 65324 13568 65340 13632
rect 65404 13568 65420 13632
rect 65484 13568 65500 13632
rect 65564 13568 65570 13632
rect 65254 13567 65570 13568
rect 64334 13088 64650 13089
rect 64334 13024 64340 13088
rect 64404 13024 64420 13088
rect 64484 13024 64500 13088
rect 64564 13024 64580 13088
rect 64644 13024 64650 13088
rect 64334 13023 64650 13024
rect 65254 12544 65570 12545
rect 65254 12480 65260 12544
rect 65324 12480 65340 12544
rect 65404 12480 65420 12544
rect 65484 12480 65500 12544
rect 65564 12480 65570 12544
rect 65254 12479 65570 12480
rect 64334 12000 64650 12001
rect 64334 11936 64340 12000
rect 64404 11936 64420 12000
rect 64484 11936 64500 12000
rect 64564 11936 64580 12000
rect 64644 11936 64650 12000
rect 64334 11935 64650 11936
rect 65254 11456 65570 11457
rect 65254 11392 65260 11456
rect 65324 11392 65340 11456
rect 65404 11392 65420 11456
rect 65484 11392 65500 11456
rect 65564 11392 65570 11456
rect 65254 11391 65570 11392
rect 64334 10912 64650 10913
rect 64334 10848 64340 10912
rect 64404 10848 64420 10912
rect 64484 10848 64500 10912
rect 64564 10848 64580 10912
rect 64644 10848 64650 10912
rect 64334 10847 64650 10848
rect 65254 10368 65570 10369
rect 65254 10304 65260 10368
rect 65324 10304 65340 10368
rect 65404 10304 65420 10368
rect 65484 10304 65500 10368
rect 65564 10304 65570 10368
rect 65254 10303 65570 10304
rect 64334 9824 64650 9825
rect 64334 9760 64340 9824
rect 64404 9760 64420 9824
rect 64484 9760 64500 9824
rect 64564 9760 64580 9824
rect 64644 9760 64650 9824
rect 64334 9759 64650 9760
rect 65254 9280 65570 9281
rect 65254 9216 65260 9280
rect 65324 9216 65340 9280
rect 65404 9216 65420 9280
rect 65484 9216 65500 9280
rect 65564 9216 65570 9280
rect 65254 9215 65570 9216
rect 64334 8736 64650 8737
rect 64334 8672 64340 8736
rect 64404 8672 64420 8736
rect 64484 8672 64500 8736
rect 64564 8672 64580 8736
rect 64644 8672 64650 8736
rect 64334 8671 64650 8672
rect 65254 8192 65570 8193
rect 65254 8128 65260 8192
rect 65324 8128 65340 8192
rect 65404 8128 65420 8192
rect 65484 8128 65500 8192
rect 65564 8128 65570 8192
rect 65254 8127 65570 8128
rect 64334 7648 64650 7649
rect 64334 7584 64340 7648
rect 64404 7584 64420 7648
rect 64484 7584 64500 7648
rect 64564 7584 64580 7648
rect 64644 7584 64650 7648
rect 64334 7583 64650 7584
rect 63534 7380 63540 7444
rect 63604 7442 63610 7444
rect 64505 7442 64571 7445
rect 63604 7440 64571 7442
rect 63604 7384 64510 7440
rect 64566 7384 64571 7440
rect 63604 7382 64571 7384
rect 63604 7380 63610 7382
rect 64505 7379 64571 7382
rect 65254 7104 65570 7105
rect 65254 7040 65260 7104
rect 65324 7040 65340 7104
rect 65404 7040 65420 7104
rect 65484 7040 65500 7104
rect 65564 7040 65570 7104
rect 65254 7039 65570 7040
rect 63902 6836 63908 6900
rect 63972 6898 63978 6900
rect 64137 6898 64203 6901
rect 64597 6898 64663 6901
rect 63972 6896 64663 6898
rect 63972 6840 64142 6896
rect 64198 6840 64602 6896
rect 64658 6840 64663 6896
rect 63972 6838 64663 6840
rect 63972 6836 63978 6838
rect 64137 6835 64203 6838
rect 64597 6835 64663 6838
rect 64334 6560 64650 6561
rect 64334 6496 64340 6560
rect 64404 6496 64420 6560
rect 64484 6496 64500 6560
rect 64564 6496 64580 6560
rect 64644 6496 64650 6560
rect 64334 6495 64650 6496
rect 65254 6016 65570 6017
rect 65254 5952 65260 6016
rect 65324 5952 65340 6016
rect 65404 5952 65420 6016
rect 65484 5952 65500 6016
rect 65564 5952 65570 6016
rect 65254 5951 65570 5952
rect 64334 5472 64650 5473
rect 64334 5408 64340 5472
rect 64404 5408 64420 5472
rect 64484 5408 64500 5472
rect 64564 5408 64580 5472
rect 64644 5408 64650 5472
rect 64334 5407 64650 5408
rect 65254 4928 65570 4929
rect 65254 4864 65260 4928
rect 65324 4864 65340 4928
rect 65404 4864 65420 4928
rect 65484 4864 65500 4928
rect 65564 4864 65570 4928
rect 65254 4863 65570 4864
rect 64334 4384 64650 4385
rect 64334 4320 64340 4384
rect 64404 4320 64420 4384
rect 64484 4320 64500 4384
rect 64564 4320 64580 4384
rect 64644 4320 64650 4384
rect 64334 4319 64650 4320
rect 65254 3840 65570 3841
rect 65254 3776 65260 3840
rect 65324 3776 65340 3840
rect 65404 3776 65420 3840
rect 65484 3776 65500 3840
rect 65564 3776 65570 3840
rect 65254 3775 65570 3776
rect 64334 3296 64650 3297
rect 64334 3232 64340 3296
rect 64404 3232 64420 3296
rect 64484 3232 64500 3296
rect 64564 3232 64580 3296
rect 64644 3232 64650 3296
rect 64334 3231 64650 3232
rect 1096 3022 1444 3044
rect 1096 2958 1118 3022
rect 1182 2958 1198 3022
rect 1262 2958 1278 3022
rect 1342 2958 1358 3022
rect 1422 2958 1444 3022
rect 1096 2942 1444 2958
rect 1096 2878 1118 2942
rect 1182 2878 1198 2942
rect 1262 2878 1278 2942
rect 1342 2878 1358 2942
rect 1422 2878 1444 2942
rect 1096 2862 1444 2878
rect 1096 2798 1118 2862
rect 1182 2798 1198 2862
rect 1262 2798 1278 2862
rect 1342 2798 1358 2862
rect 1422 2798 1444 2862
rect 1096 2782 1444 2798
rect 1096 2718 1118 2782
rect 1182 2718 1198 2782
rect 1262 2718 1278 2782
rect 1342 2718 1358 2782
rect 1422 2718 1444 2782
rect 1096 2696 1444 2718
rect 61492 3022 61840 3044
rect 61492 2958 61514 3022
rect 61578 2958 61594 3022
rect 61658 2958 61674 3022
rect 61738 2958 61754 3022
rect 61818 2958 61840 3022
rect 61492 2942 61840 2958
rect 61492 2878 61514 2942
rect 61578 2878 61594 2942
rect 61658 2878 61674 2942
rect 61738 2878 61754 2942
rect 61818 2878 61840 2942
rect 61492 2862 61840 2878
rect 61492 2798 61514 2862
rect 61578 2798 61594 2862
rect 61658 2798 61674 2862
rect 61738 2798 61754 2862
rect 61818 2798 61840 2862
rect 61492 2782 61840 2798
rect 61492 2718 61514 2782
rect 61578 2718 61594 2782
rect 61658 2718 61674 2782
rect 61738 2718 61754 2782
rect 61818 2718 61840 2782
rect 61492 2696 61840 2718
rect 65254 2752 65570 2753
rect 65254 2688 65260 2752
rect 65324 2688 65340 2752
rect 65404 2688 65420 2752
rect 65484 2688 65500 2752
rect 65564 2688 65570 2752
rect 65254 2687 65570 2688
rect 400 2326 748 2348
rect 400 2262 422 2326
rect 486 2262 502 2326
rect 566 2262 582 2326
rect 646 2262 662 2326
rect 726 2262 748 2326
rect 400 2246 748 2262
rect 400 2182 422 2246
rect 486 2182 502 2246
rect 566 2182 582 2246
rect 646 2182 662 2246
rect 726 2182 748 2246
rect 400 2166 748 2182
rect 400 2102 422 2166
rect 486 2102 502 2166
rect 566 2102 582 2166
rect 646 2102 662 2166
rect 726 2102 748 2166
rect 400 2086 748 2102
rect 400 2022 422 2086
rect 486 2022 502 2086
rect 566 2022 582 2086
rect 646 2022 662 2086
rect 726 2022 748 2086
rect 400 2000 748 2022
rect 62188 2326 62536 2348
rect 62188 2262 62210 2326
rect 62274 2262 62290 2326
rect 62354 2262 62370 2326
rect 62434 2262 62450 2326
rect 62514 2262 62536 2326
rect 62188 2246 62536 2262
rect 62188 2182 62210 2246
rect 62274 2182 62290 2246
rect 62354 2182 62370 2246
rect 62434 2182 62450 2246
rect 62514 2182 62536 2246
rect 62188 2166 62536 2182
rect 62188 2102 62210 2166
rect 62274 2102 62290 2166
rect 62354 2102 62370 2166
rect 62434 2102 62450 2166
rect 62514 2102 62536 2166
rect 64334 2208 64650 2209
rect 64334 2144 64340 2208
rect 64404 2144 64420 2208
rect 64484 2144 64500 2208
rect 64564 2144 64580 2208
rect 64644 2144 64650 2208
rect 64334 2143 64650 2144
rect 62188 2086 62536 2102
rect 62188 2022 62210 2086
rect 62274 2022 62290 2086
rect 62354 2022 62370 2086
rect 62434 2022 62450 2086
rect 62514 2022 62536 2086
rect 62188 2000 62536 2022
rect 48957 1868 49023 1869
rect 48935 1866 48941 1868
rect 48866 1806 48941 1866
rect 49005 1864 49023 1868
rect 49018 1808 49023 1864
rect 48935 1804 48941 1806
rect 49005 1804 49023 1808
rect 49366 1804 49372 1868
rect 49436 1866 49442 1868
rect 49601 1866 49667 1869
rect 63677 1866 63743 1869
rect 49436 1864 49667 1866
rect 49436 1808 49606 1864
rect 49662 1808 49667 1864
rect 49436 1806 49667 1808
rect 49436 1804 49442 1806
rect 48957 1803 49023 1804
rect 49601 1803 49667 1806
rect 55170 1864 63743 1866
rect 55170 1808 63682 1864
rect 63738 1808 63743 1864
rect 55170 1806 63743 1808
rect 49693 1732 49759 1733
rect 49668 1730 49674 1732
rect 49602 1670 49674 1730
rect 49738 1728 49759 1732
rect 49754 1672 49759 1728
rect 49668 1668 49674 1670
rect 49738 1668 49759 1672
rect 49693 1667 49759 1668
rect 49073 1532 49079 1596
rect 49143 1532 49149 1596
rect 49211 1532 49217 1596
rect 49281 1594 49287 1596
rect 55170 1594 55230 1806
rect 63677 1803 63743 1806
rect 65254 1664 65570 1665
rect 65254 1600 65260 1664
rect 65324 1600 65340 1664
rect 65404 1600 65420 1664
rect 65484 1600 65500 1664
rect 65564 1600 65570 1664
rect 65254 1599 65570 1600
rect 49281 1534 55230 1594
rect 49281 1532 49287 1534
rect 49081 1458 49141 1532
rect 62757 1458 62823 1461
rect 49081 1456 62823 1458
rect 49081 1400 62762 1456
rect 62818 1400 62823 1456
rect 49081 1398 62823 1400
rect 62757 1395 62823 1398
rect 49918 1260 49924 1324
rect 49988 1322 49994 1324
rect 62941 1322 63007 1325
rect 49988 1320 63007 1322
rect 49988 1264 62946 1320
rect 63002 1264 63007 1320
rect 49988 1262 63007 1264
rect 49988 1260 49994 1262
rect 62941 1259 63007 1262
rect 64334 1120 64650 1121
rect 64334 1056 64340 1120
rect 64404 1056 64420 1120
rect 64484 1056 64500 1120
rect 64564 1056 64580 1120
rect 64644 1056 64650 1120
rect 64334 1055 64650 1056
rect 65254 576 65570 577
rect 65254 512 65260 576
rect 65324 512 65340 576
rect 65404 512 65420 576
rect 65484 512 65500 576
rect 65564 512 65570 576
rect 65254 511 65570 512
<< via3 >>
rect 26004 44916 26068 44980
rect 13308 44780 13372 44844
rect 13860 44840 13924 44844
rect 13860 44784 13874 44840
rect 13874 44784 13924 44840
rect 13860 44780 13924 44784
rect 27660 44780 27724 44844
rect 11652 44644 11716 44708
rect 14964 44644 15028 44708
rect 27108 44644 27172 44708
rect 28212 44644 28276 44708
rect 2000 44636 2064 44640
rect 2000 44580 2004 44636
rect 2004 44580 2060 44636
rect 2060 44580 2064 44636
rect 2000 44576 2064 44580
rect 2080 44636 2144 44640
rect 2080 44580 2084 44636
rect 2084 44580 2140 44636
rect 2140 44580 2144 44636
rect 2080 44576 2144 44580
rect 2160 44636 2224 44640
rect 2160 44580 2164 44636
rect 2164 44580 2220 44636
rect 2220 44580 2224 44636
rect 2160 44576 2224 44580
rect 2240 44636 2304 44640
rect 2240 44580 2244 44636
rect 2244 44580 2300 44636
rect 2300 44580 2304 44636
rect 2240 44576 2304 44580
rect 50000 44636 50064 44640
rect 50000 44580 50004 44636
rect 50004 44580 50060 44636
rect 50060 44580 50064 44636
rect 50000 44576 50064 44580
rect 50080 44636 50144 44640
rect 50080 44580 50084 44636
rect 50084 44580 50140 44636
rect 50140 44580 50144 44636
rect 50080 44576 50144 44580
rect 50160 44636 50224 44640
rect 50160 44580 50164 44636
rect 50164 44580 50220 44636
rect 50220 44580 50224 44636
rect 50160 44576 50224 44580
rect 50240 44636 50304 44640
rect 50240 44580 50244 44636
rect 50244 44580 50300 44636
rect 50300 44580 50304 44636
rect 50240 44576 50304 44580
rect 6132 44568 6196 44572
rect 6132 44512 6182 44568
rect 6182 44512 6196 44568
rect 6132 44508 6196 44512
rect 6684 44568 6748 44572
rect 6684 44512 6734 44568
rect 6734 44512 6748 44568
rect 6684 44508 6748 44512
rect 7236 44568 7300 44572
rect 7236 44512 7286 44568
rect 7286 44512 7300 44568
rect 7236 44508 7300 44512
rect 7788 44568 7852 44572
rect 7788 44512 7838 44568
rect 7838 44512 7852 44568
rect 7788 44508 7852 44512
rect 8340 44568 8404 44572
rect 8340 44512 8390 44568
rect 8390 44512 8404 44568
rect 8340 44508 8404 44512
rect 8892 44568 8956 44572
rect 8892 44512 8942 44568
rect 8942 44512 8956 44568
rect 8892 44508 8956 44512
rect 9444 44568 9508 44572
rect 9444 44512 9494 44568
rect 9494 44512 9508 44568
rect 9444 44508 9508 44512
rect 9996 44568 10060 44572
rect 9996 44512 10046 44568
rect 10046 44512 10060 44568
rect 9996 44508 10060 44512
rect 10548 44568 10612 44572
rect 10548 44512 10562 44568
rect 10562 44512 10612 44568
rect 10548 44508 10612 44512
rect 11100 44508 11164 44572
rect 12204 44508 12268 44572
rect 14412 44508 14476 44572
rect 15516 44508 15580 44572
rect 17724 44508 17788 44572
rect 26556 44372 26620 44436
rect 2920 44092 2984 44096
rect 2920 44036 2924 44092
rect 2924 44036 2980 44092
rect 2980 44036 2984 44092
rect 2920 44032 2984 44036
rect 3000 44092 3064 44096
rect 3000 44036 3004 44092
rect 3004 44036 3060 44092
rect 3060 44036 3064 44092
rect 3000 44032 3064 44036
rect 3080 44092 3144 44096
rect 3080 44036 3084 44092
rect 3084 44036 3140 44092
rect 3140 44036 3144 44092
rect 3080 44032 3144 44036
rect 3160 44092 3224 44096
rect 3160 44036 3164 44092
rect 3164 44036 3220 44092
rect 3220 44036 3224 44092
rect 3160 44032 3224 44036
rect 50920 44092 50984 44096
rect 50920 44036 50924 44092
rect 50924 44036 50980 44092
rect 50980 44036 50984 44092
rect 50920 44032 50984 44036
rect 51000 44092 51064 44096
rect 51000 44036 51004 44092
rect 51004 44036 51060 44092
rect 51060 44036 51064 44092
rect 51000 44032 51064 44036
rect 51080 44092 51144 44096
rect 51080 44036 51084 44092
rect 51084 44036 51140 44092
rect 51140 44036 51144 44092
rect 51080 44032 51144 44036
rect 51160 44092 51224 44096
rect 51160 44036 51164 44092
rect 51164 44036 51220 44092
rect 51220 44036 51224 44092
rect 51160 44032 51224 44036
rect 18276 44024 18340 44028
rect 18276 43968 18326 44024
rect 18326 43968 18340 44024
rect 18276 43964 18340 43968
rect 12756 43888 12820 43892
rect 12756 43832 12806 43888
rect 12806 43832 12820 43888
rect 12756 43828 12820 43832
rect 16068 43828 16132 43892
rect 2000 43548 2064 43552
rect 2000 43492 2004 43548
rect 2004 43492 2060 43548
rect 2060 43492 2064 43548
rect 2000 43488 2064 43492
rect 2080 43548 2144 43552
rect 2080 43492 2084 43548
rect 2084 43492 2140 43548
rect 2140 43492 2144 43548
rect 2080 43488 2144 43492
rect 2160 43548 2224 43552
rect 2160 43492 2164 43548
rect 2164 43492 2220 43548
rect 2220 43492 2224 43548
rect 2160 43488 2224 43492
rect 2240 43548 2304 43552
rect 2240 43492 2244 43548
rect 2244 43492 2300 43548
rect 2300 43492 2304 43548
rect 2240 43488 2304 43492
rect 17172 43420 17236 43484
rect 23244 43420 23308 43484
rect 50000 43548 50064 43552
rect 50000 43492 50004 43548
rect 50004 43492 50060 43548
rect 50060 43492 50064 43548
rect 50000 43488 50064 43492
rect 50080 43548 50144 43552
rect 50080 43492 50084 43548
rect 50084 43492 50140 43548
rect 50140 43492 50144 43548
rect 50080 43488 50144 43492
rect 50160 43548 50224 43552
rect 50160 43492 50164 43548
rect 50164 43492 50220 43548
rect 50220 43492 50224 43548
rect 50160 43488 50224 43492
rect 50240 43548 50304 43552
rect 50240 43492 50244 43548
rect 50244 43492 50300 43548
rect 50300 43492 50304 43548
rect 50240 43488 50304 43492
rect 22140 43284 22204 43348
rect 24716 43284 24780 43348
rect 32076 43420 32140 43484
rect 35204 43148 35268 43212
rect 27476 43012 27540 43076
rect 27660 43012 27724 43076
rect 2920 43004 2984 43008
rect 2920 42948 2924 43004
rect 2924 42948 2980 43004
rect 2980 42948 2984 43004
rect 2920 42944 2984 42948
rect 3000 43004 3064 43008
rect 3000 42948 3004 43004
rect 3004 42948 3060 43004
rect 3060 42948 3064 43004
rect 3000 42944 3064 42948
rect 3080 43004 3144 43008
rect 3080 42948 3084 43004
rect 3084 42948 3140 43004
rect 3140 42948 3144 43004
rect 3080 42944 3144 42948
rect 3160 43004 3224 43008
rect 3160 42948 3164 43004
rect 3164 42948 3220 43004
rect 3220 42948 3224 43004
rect 3160 42944 3224 42948
rect 50920 43004 50984 43008
rect 50920 42948 50924 43004
rect 50924 42948 50980 43004
rect 50980 42948 50984 43004
rect 50920 42944 50984 42948
rect 51000 43004 51064 43008
rect 51000 42948 51004 43004
rect 51004 42948 51060 43004
rect 51060 42948 51064 43004
rect 51000 42944 51064 42948
rect 51080 43004 51144 43008
rect 51080 42948 51084 43004
rect 51084 42948 51140 43004
rect 51140 42948 51144 43004
rect 51080 42944 51144 42948
rect 51160 43004 51224 43008
rect 51160 42948 51164 43004
rect 51164 42948 51220 43004
rect 51220 42948 51224 43004
rect 51160 42944 51224 42948
rect 16620 42876 16684 42940
rect 24900 42876 24964 42940
rect 2000 42460 2064 42464
rect 2000 42404 2004 42460
rect 2004 42404 2060 42460
rect 2060 42404 2064 42460
rect 2000 42400 2064 42404
rect 2080 42460 2144 42464
rect 2080 42404 2084 42460
rect 2084 42404 2140 42460
rect 2140 42404 2144 42460
rect 2080 42400 2144 42404
rect 2160 42460 2224 42464
rect 2160 42404 2164 42460
rect 2164 42404 2220 42460
rect 2220 42404 2224 42460
rect 2160 42400 2224 42404
rect 2240 42460 2304 42464
rect 2240 42404 2244 42460
rect 2244 42404 2300 42460
rect 2300 42404 2304 42460
rect 2240 42400 2304 42404
rect 50000 42460 50064 42464
rect 50000 42404 50004 42460
rect 50004 42404 50060 42460
rect 50060 42404 50064 42460
rect 50000 42400 50064 42404
rect 50080 42460 50144 42464
rect 50080 42404 50084 42460
rect 50084 42404 50140 42460
rect 50140 42404 50144 42460
rect 50080 42400 50144 42404
rect 50160 42460 50224 42464
rect 50160 42404 50164 42460
rect 50164 42404 50220 42460
rect 50220 42404 50224 42460
rect 50160 42400 50224 42404
rect 50240 42460 50304 42464
rect 50240 42404 50244 42460
rect 50244 42404 50300 42460
rect 50300 42404 50304 42460
rect 50240 42400 50304 42404
rect 18828 42332 18892 42396
rect 30972 42060 31036 42124
rect 2920 41916 2984 41920
rect 2920 41860 2924 41916
rect 2924 41860 2980 41916
rect 2980 41860 2984 41916
rect 2920 41856 2984 41860
rect 3000 41916 3064 41920
rect 3000 41860 3004 41916
rect 3004 41860 3060 41916
rect 3060 41860 3064 41916
rect 3000 41856 3064 41860
rect 3080 41916 3144 41920
rect 3080 41860 3084 41916
rect 3084 41860 3140 41916
rect 3140 41860 3144 41916
rect 3080 41856 3144 41860
rect 3160 41916 3224 41920
rect 3160 41860 3164 41916
rect 3164 41860 3220 41916
rect 3220 41860 3224 41916
rect 3160 41856 3224 41860
rect 50920 41916 50984 41920
rect 50920 41860 50924 41916
rect 50924 41860 50980 41916
rect 50980 41860 50984 41916
rect 50920 41856 50984 41860
rect 51000 41916 51064 41920
rect 51000 41860 51004 41916
rect 51004 41860 51060 41916
rect 51060 41860 51064 41916
rect 51000 41856 51064 41860
rect 51080 41916 51144 41920
rect 51080 41860 51084 41916
rect 51084 41860 51140 41916
rect 51140 41860 51144 41916
rect 51080 41856 51144 41860
rect 51160 41916 51224 41920
rect 51160 41860 51164 41916
rect 51164 41860 51220 41916
rect 51220 41860 51224 41916
rect 51160 41856 51224 41860
rect 2000 41372 2064 41376
rect 2000 41316 2004 41372
rect 2004 41316 2060 41372
rect 2060 41316 2064 41372
rect 2000 41312 2064 41316
rect 2080 41372 2144 41376
rect 2080 41316 2084 41372
rect 2084 41316 2140 41372
rect 2140 41316 2144 41372
rect 2080 41312 2144 41316
rect 2160 41372 2224 41376
rect 2160 41316 2164 41372
rect 2164 41316 2220 41372
rect 2220 41316 2224 41372
rect 2160 41312 2224 41316
rect 2240 41372 2304 41376
rect 2240 41316 2244 41372
rect 2244 41316 2300 41372
rect 2300 41316 2304 41372
rect 2240 41312 2304 41316
rect 50000 41372 50064 41376
rect 50000 41316 50004 41372
rect 50004 41316 50060 41372
rect 50060 41316 50064 41372
rect 50000 41312 50064 41316
rect 50080 41372 50144 41376
rect 50080 41316 50084 41372
rect 50084 41316 50140 41372
rect 50140 41316 50144 41372
rect 50080 41312 50144 41316
rect 50160 41372 50224 41376
rect 50160 41316 50164 41372
rect 50164 41316 50220 41372
rect 50220 41316 50224 41372
rect 50160 41312 50224 41316
rect 50240 41372 50304 41376
rect 50240 41316 50244 41372
rect 50244 41316 50300 41372
rect 50300 41316 50304 41372
rect 50240 41312 50304 41316
rect 35020 41244 35084 41308
rect 26924 40972 26988 41036
rect 32996 40836 33060 40900
rect 2920 40828 2984 40832
rect 2920 40772 2924 40828
rect 2924 40772 2980 40828
rect 2980 40772 2984 40828
rect 2920 40768 2984 40772
rect 3000 40828 3064 40832
rect 3000 40772 3004 40828
rect 3004 40772 3060 40828
rect 3060 40772 3064 40828
rect 3000 40768 3064 40772
rect 3080 40828 3144 40832
rect 3080 40772 3084 40828
rect 3084 40772 3140 40828
rect 3140 40772 3144 40828
rect 3080 40768 3144 40772
rect 3160 40828 3224 40832
rect 3160 40772 3164 40828
rect 3164 40772 3220 40828
rect 3220 40772 3224 40828
rect 3160 40768 3224 40772
rect 50920 40828 50984 40832
rect 50920 40772 50924 40828
rect 50924 40772 50980 40828
rect 50980 40772 50984 40828
rect 50920 40768 50984 40772
rect 51000 40828 51064 40832
rect 51000 40772 51004 40828
rect 51004 40772 51060 40828
rect 51060 40772 51064 40828
rect 51000 40768 51064 40772
rect 51080 40828 51144 40832
rect 51080 40772 51084 40828
rect 51084 40772 51140 40828
rect 51140 40772 51144 40828
rect 51080 40768 51144 40772
rect 51160 40828 51224 40832
rect 51160 40772 51164 40828
rect 51164 40772 51220 40828
rect 51220 40772 51224 40828
rect 51160 40768 51224 40772
rect 27476 40700 27540 40764
rect 3924 40564 3988 40628
rect 23796 40564 23860 40628
rect 25452 40564 25516 40628
rect 32812 40564 32876 40628
rect 27844 40292 27908 40356
rect 2000 40284 2064 40288
rect 2000 40228 2004 40284
rect 2004 40228 2060 40284
rect 2060 40228 2064 40284
rect 2000 40224 2064 40228
rect 2080 40284 2144 40288
rect 2080 40228 2084 40284
rect 2084 40228 2140 40284
rect 2140 40228 2144 40284
rect 2080 40224 2144 40228
rect 2160 40284 2224 40288
rect 2160 40228 2164 40284
rect 2164 40228 2220 40284
rect 2220 40228 2224 40284
rect 2160 40224 2224 40228
rect 2240 40284 2304 40288
rect 2240 40228 2244 40284
rect 2244 40228 2300 40284
rect 2300 40228 2304 40284
rect 2240 40224 2304 40228
rect 50000 40284 50064 40288
rect 50000 40228 50004 40284
rect 50004 40228 50060 40284
rect 50060 40228 50064 40284
rect 50000 40224 50064 40228
rect 50080 40284 50144 40288
rect 50080 40228 50084 40284
rect 50084 40228 50140 40284
rect 50140 40228 50144 40284
rect 50080 40224 50144 40228
rect 50160 40284 50224 40288
rect 50160 40228 50164 40284
rect 50164 40228 50220 40284
rect 50220 40228 50224 40284
rect 50160 40224 50224 40228
rect 50240 40284 50304 40288
rect 50240 40228 50244 40284
rect 50244 40228 50300 40284
rect 50300 40228 50304 40284
rect 50240 40224 50304 40228
rect 24348 40020 24412 40084
rect 28580 39884 28644 39948
rect 15516 39748 15580 39812
rect 2920 39740 2984 39744
rect 2920 39684 2924 39740
rect 2924 39684 2980 39740
rect 2980 39684 2984 39740
rect 2920 39680 2984 39684
rect 3000 39740 3064 39744
rect 3000 39684 3004 39740
rect 3004 39684 3060 39740
rect 3060 39684 3064 39740
rect 3000 39680 3064 39684
rect 3080 39740 3144 39744
rect 3080 39684 3084 39740
rect 3084 39684 3140 39740
rect 3140 39684 3144 39740
rect 3080 39680 3144 39684
rect 3160 39740 3224 39744
rect 3160 39684 3164 39740
rect 3164 39684 3220 39740
rect 3220 39684 3224 39740
rect 3160 39680 3224 39684
rect 50920 39740 50984 39744
rect 50920 39684 50924 39740
rect 50924 39684 50980 39740
rect 50980 39684 50984 39740
rect 50920 39680 50984 39684
rect 51000 39740 51064 39744
rect 51000 39684 51004 39740
rect 51004 39684 51060 39740
rect 51060 39684 51064 39740
rect 51000 39680 51064 39684
rect 51080 39740 51144 39744
rect 51080 39684 51084 39740
rect 51084 39684 51140 39740
rect 51140 39684 51144 39740
rect 51080 39680 51144 39684
rect 51160 39740 51224 39744
rect 51160 39684 51164 39740
rect 51164 39684 51220 39740
rect 51220 39684 51224 39740
rect 51160 39680 51224 39684
rect 32996 39612 33060 39676
rect 36124 39612 36188 39676
rect 19012 39340 19076 39404
rect 27844 39204 27908 39268
rect 32812 39204 32876 39268
rect 2000 39196 2064 39200
rect 2000 39140 2004 39196
rect 2004 39140 2060 39196
rect 2060 39140 2064 39196
rect 2000 39136 2064 39140
rect 2080 39196 2144 39200
rect 2080 39140 2084 39196
rect 2084 39140 2140 39196
rect 2140 39140 2144 39196
rect 2080 39136 2144 39140
rect 2160 39196 2224 39200
rect 2160 39140 2164 39196
rect 2164 39140 2220 39196
rect 2220 39140 2224 39196
rect 2160 39136 2224 39140
rect 2240 39196 2304 39200
rect 2240 39140 2244 39196
rect 2244 39140 2300 39196
rect 2300 39140 2304 39196
rect 2240 39136 2304 39140
rect 50000 39196 50064 39200
rect 50000 39140 50004 39196
rect 50004 39140 50060 39196
rect 50060 39140 50064 39196
rect 50000 39136 50064 39140
rect 50080 39196 50144 39200
rect 50080 39140 50084 39196
rect 50084 39140 50140 39196
rect 50140 39140 50144 39196
rect 50080 39136 50144 39140
rect 50160 39196 50224 39200
rect 50160 39140 50164 39196
rect 50164 39140 50220 39196
rect 50220 39140 50224 39196
rect 50160 39136 50224 39140
rect 50240 39196 50304 39200
rect 50240 39140 50244 39196
rect 50244 39140 50300 39196
rect 50300 39140 50304 39196
rect 50240 39136 50304 39140
rect 28948 38932 29012 38996
rect 26188 38660 26252 38724
rect 28396 38660 28460 38724
rect 32444 38660 32508 38724
rect 2920 38652 2984 38656
rect 2920 38596 2924 38652
rect 2924 38596 2980 38652
rect 2980 38596 2984 38652
rect 2920 38592 2984 38596
rect 3000 38652 3064 38656
rect 3000 38596 3004 38652
rect 3004 38596 3060 38652
rect 3060 38596 3064 38652
rect 3000 38592 3064 38596
rect 3080 38652 3144 38656
rect 3080 38596 3084 38652
rect 3084 38596 3140 38652
rect 3140 38596 3144 38652
rect 3080 38592 3144 38596
rect 3160 38652 3224 38656
rect 3160 38596 3164 38652
rect 3164 38596 3220 38652
rect 3220 38596 3224 38652
rect 3160 38592 3224 38596
rect 24532 38584 24596 38588
rect 24532 38528 24582 38584
rect 24582 38528 24596 38584
rect 24532 38524 24596 38528
rect 33180 38660 33244 38724
rect 35388 38660 35452 38724
rect 46980 38660 47044 38724
rect 50920 38652 50984 38656
rect 50920 38596 50924 38652
rect 50924 38596 50980 38652
rect 50980 38596 50984 38652
rect 50920 38592 50984 38596
rect 51000 38652 51064 38656
rect 51000 38596 51004 38652
rect 51004 38596 51060 38652
rect 51060 38596 51064 38652
rect 51000 38592 51064 38596
rect 51080 38652 51144 38656
rect 51080 38596 51084 38652
rect 51084 38596 51140 38652
rect 51140 38596 51144 38652
rect 51080 38592 51144 38596
rect 51160 38652 51224 38656
rect 51160 38596 51164 38652
rect 51164 38596 51220 38652
rect 51220 38596 51224 38652
rect 51160 38592 51224 38596
rect 26004 38388 26068 38452
rect 34100 38524 34164 38588
rect 62804 38524 62868 38588
rect 21404 38252 21468 38316
rect 2000 38108 2064 38112
rect 2000 38052 2004 38108
rect 2004 38052 2060 38108
rect 2060 38052 2064 38108
rect 2000 38048 2064 38052
rect 2080 38108 2144 38112
rect 2080 38052 2084 38108
rect 2084 38052 2140 38108
rect 2140 38052 2144 38108
rect 2080 38048 2144 38052
rect 2160 38108 2224 38112
rect 2160 38052 2164 38108
rect 2164 38052 2220 38108
rect 2220 38052 2224 38108
rect 2160 38048 2224 38052
rect 2240 38108 2304 38112
rect 2240 38052 2244 38108
rect 2244 38052 2300 38108
rect 2300 38052 2304 38108
rect 2240 38048 2304 38052
rect 20116 37980 20180 38044
rect 28028 37844 28092 37908
rect 50000 38108 50064 38112
rect 50000 38052 50004 38108
rect 50004 38052 50060 38108
rect 50060 38052 50064 38108
rect 50000 38048 50064 38052
rect 50080 38108 50144 38112
rect 50080 38052 50084 38108
rect 50084 38052 50140 38108
rect 50140 38052 50144 38108
rect 50080 38048 50144 38052
rect 50160 38108 50224 38112
rect 50160 38052 50164 38108
rect 50164 38052 50220 38108
rect 50220 38052 50224 38108
rect 50160 38048 50224 38052
rect 50240 38108 50304 38112
rect 50240 38052 50244 38108
rect 50244 38052 50300 38108
rect 50300 38052 50304 38108
rect 50240 38048 50304 38052
rect 62988 37708 63052 37772
rect 2920 37564 2984 37568
rect 2920 37508 2924 37564
rect 2924 37508 2980 37564
rect 2980 37508 2984 37564
rect 2920 37504 2984 37508
rect 3000 37564 3064 37568
rect 3000 37508 3004 37564
rect 3004 37508 3060 37564
rect 3060 37508 3064 37564
rect 3000 37504 3064 37508
rect 3080 37564 3144 37568
rect 3080 37508 3084 37564
rect 3084 37508 3140 37564
rect 3140 37508 3144 37564
rect 3080 37504 3144 37508
rect 3160 37564 3224 37568
rect 3160 37508 3164 37564
rect 3164 37508 3220 37564
rect 3220 37508 3224 37564
rect 3160 37504 3224 37508
rect 50920 37564 50984 37568
rect 50920 37508 50924 37564
rect 50924 37508 50980 37564
rect 50980 37508 50984 37564
rect 50920 37504 50984 37508
rect 51000 37564 51064 37568
rect 51000 37508 51004 37564
rect 51004 37508 51060 37564
rect 51060 37508 51064 37564
rect 51000 37504 51064 37508
rect 51080 37564 51144 37568
rect 51080 37508 51084 37564
rect 51084 37508 51140 37564
rect 51140 37508 51144 37564
rect 51080 37504 51144 37508
rect 51160 37564 51224 37568
rect 51160 37508 51164 37564
rect 51164 37508 51220 37564
rect 51220 37508 51224 37564
rect 51160 37504 51224 37508
rect 65260 37564 65324 37568
rect 65260 37508 65264 37564
rect 65264 37508 65320 37564
rect 65320 37508 65324 37564
rect 65260 37504 65324 37508
rect 65340 37564 65404 37568
rect 65340 37508 65344 37564
rect 65344 37508 65400 37564
rect 65400 37508 65404 37564
rect 65340 37504 65404 37508
rect 65420 37564 65484 37568
rect 65420 37508 65424 37564
rect 65424 37508 65480 37564
rect 65480 37508 65484 37564
rect 65420 37504 65484 37508
rect 65500 37564 65564 37568
rect 65500 37508 65504 37564
rect 65504 37508 65560 37564
rect 65560 37508 65564 37564
rect 65500 37504 65564 37508
rect 27292 37436 27356 37500
rect 28580 37496 28644 37500
rect 28580 37440 28594 37496
rect 28594 37440 28644 37496
rect 28580 37436 28644 37440
rect 31892 37436 31956 37500
rect 32996 37436 33060 37500
rect 24716 37300 24780 37364
rect 27844 37300 27908 37364
rect 14412 37164 14476 37228
rect 22692 37164 22756 37228
rect 24900 37164 24964 37228
rect 28212 37164 28276 37228
rect 45876 37300 45940 37364
rect 12020 37028 12084 37092
rect 23612 37028 23676 37092
rect 2000 37020 2064 37024
rect 2000 36964 2004 37020
rect 2004 36964 2060 37020
rect 2060 36964 2064 37020
rect 2000 36960 2064 36964
rect 2080 37020 2144 37024
rect 2080 36964 2084 37020
rect 2084 36964 2140 37020
rect 2140 36964 2144 37020
rect 2080 36960 2144 36964
rect 2160 37020 2224 37024
rect 2160 36964 2164 37020
rect 2164 36964 2220 37020
rect 2220 36964 2224 37020
rect 2160 36960 2224 36964
rect 2240 37020 2304 37024
rect 2240 36964 2244 37020
rect 2244 36964 2300 37020
rect 2300 36964 2304 37020
rect 2240 36960 2304 36964
rect 50000 37020 50064 37024
rect 50000 36964 50004 37020
rect 50004 36964 50060 37020
rect 50060 36964 50064 37020
rect 50000 36960 50064 36964
rect 50080 37020 50144 37024
rect 50080 36964 50084 37020
rect 50084 36964 50140 37020
rect 50140 36964 50144 37020
rect 50080 36960 50144 36964
rect 50160 37020 50224 37024
rect 50160 36964 50164 37020
rect 50164 36964 50220 37020
rect 50220 36964 50224 37020
rect 50160 36960 50224 36964
rect 50240 37020 50304 37024
rect 50240 36964 50244 37020
rect 50244 36964 50300 37020
rect 50300 36964 50304 37020
rect 50240 36960 50304 36964
rect 64340 37020 64404 37024
rect 64340 36964 64344 37020
rect 64344 36964 64400 37020
rect 64400 36964 64404 37020
rect 64340 36960 64404 36964
rect 64420 37020 64484 37024
rect 64420 36964 64424 37020
rect 64424 36964 64480 37020
rect 64480 36964 64484 37020
rect 64420 36960 64484 36964
rect 64500 37020 64564 37024
rect 64500 36964 64504 37020
rect 64504 36964 64560 37020
rect 64560 36964 64564 37020
rect 64500 36960 64564 36964
rect 64580 37020 64644 37024
rect 64580 36964 64584 37020
rect 64584 36964 64640 37020
rect 64640 36964 64644 37020
rect 64580 36960 64644 36964
rect 10916 36892 10980 36956
rect 38884 36892 38948 36956
rect 9628 36756 9692 36820
rect 37596 36756 37660 36820
rect 62620 36756 62684 36820
rect 5028 36620 5092 36684
rect 39988 36620 40052 36684
rect 6132 36484 6196 36548
rect 26740 36484 26804 36548
rect 65260 36476 65324 36480
rect 65260 36420 65264 36476
rect 65264 36420 65320 36476
rect 65320 36420 65324 36476
rect 65260 36416 65324 36420
rect 65340 36476 65404 36480
rect 65340 36420 65344 36476
rect 65344 36420 65400 36476
rect 65400 36420 65404 36476
rect 65340 36416 65404 36420
rect 65420 36476 65484 36480
rect 65420 36420 65424 36476
rect 65424 36420 65480 36476
rect 65480 36420 65484 36476
rect 65420 36416 65484 36420
rect 65500 36476 65564 36480
rect 65500 36420 65504 36476
rect 65504 36420 65560 36476
rect 65560 36420 65564 36476
rect 65500 36416 65564 36420
rect 22508 36348 22572 36412
rect 33180 36348 33244 36412
rect 21588 36212 21652 36276
rect 16620 36076 16684 36140
rect 13158 35940 13222 36004
rect 17830 35804 17894 35868
rect 19472 35804 19536 35868
rect 20968 35804 21032 35868
rect 23198 35864 23262 35868
rect 23198 35808 23202 35864
rect 23202 35808 23258 35864
rect 23258 35808 23262 35864
rect 23198 35804 23262 35808
rect 24692 36000 24756 36004
rect 24692 35944 24730 36000
rect 24730 35944 24756 36000
rect 24692 35940 24756 35944
rect 26464 35940 26528 36004
rect 29198 35940 29262 36004
rect 30678 36000 30742 36004
rect 30678 35944 30710 36000
rect 30710 35944 30742 36000
rect 25868 35864 25932 35868
rect 25868 35808 25870 35864
rect 25870 35808 25926 35864
rect 25926 35808 25932 35864
rect 25868 35804 25932 35808
rect 29510 35804 29574 35868
rect 30236 35864 30300 35868
rect 30236 35808 30286 35864
rect 30286 35808 30300 35864
rect 30236 35804 30300 35808
rect 30678 35940 30742 35944
rect 31198 35940 31262 36004
rect 31708 35940 31772 36004
rect 32076 35940 32140 36004
rect 33916 35804 33980 35868
rect 36518 35804 36582 35868
rect 42358 35804 42422 35868
rect 43526 35864 43590 35868
rect 43526 35808 43534 35864
rect 43534 35808 43590 35864
rect 43526 35804 43590 35808
rect 64092 35940 64156 36004
rect 64340 35932 64404 35936
rect 64340 35876 64344 35932
rect 64344 35876 64400 35932
rect 64400 35876 64404 35932
rect 64340 35872 64404 35876
rect 64420 35932 64484 35936
rect 64420 35876 64424 35932
rect 64424 35876 64480 35932
rect 64480 35876 64484 35932
rect 64420 35872 64484 35876
rect 64500 35932 64564 35936
rect 64500 35876 64504 35932
rect 64504 35876 64560 35932
rect 64560 35876 64564 35932
rect 64500 35872 64564 35876
rect 64580 35932 64644 35936
rect 64580 35876 64584 35932
rect 64584 35876 64640 35932
rect 64640 35876 64644 35932
rect 64580 35872 64644 35876
rect 63540 35804 63604 35868
rect 7328 35668 7392 35732
rect 8486 35728 8550 35732
rect 8486 35672 8538 35728
rect 8538 35672 8550 35728
rect 8486 35668 8550 35672
rect 20028 35728 20092 35732
rect 20028 35672 20074 35728
rect 20074 35672 20092 35728
rect 20028 35668 20092 35672
rect 21196 35728 21260 35732
rect 21196 35672 21234 35728
rect 21234 35672 21260 35728
rect 21196 35668 21260 35672
rect 21968 35728 22032 35732
rect 21968 35672 22006 35728
rect 22006 35672 22032 35728
rect 21968 35668 22032 35672
rect 22140 35728 22204 35732
rect 22140 35672 22190 35728
rect 22190 35672 22204 35728
rect 22140 35668 22204 35672
rect 22968 35728 23032 35732
rect 22968 35672 23018 35728
rect 23018 35672 23032 35728
rect 22968 35668 23032 35672
rect 23532 35728 23596 35732
rect 23532 35672 23570 35728
rect 23570 35672 23596 35728
rect 23532 35668 23596 35672
rect 25210 35668 25274 35732
rect 26188 35668 26252 35732
rect 29968 35728 30032 35732
rect 29968 35672 30010 35728
rect 30010 35672 30032 35728
rect 29968 35668 30032 35672
rect 32876 35668 32940 35732
rect 33456 35668 33520 35732
rect 33732 35668 33796 35732
rect 41184 35668 41248 35732
rect 44680 35668 44744 35732
rect 56246 35668 56310 35732
rect 62804 35532 62868 35596
rect 422 35428 486 35492
rect 502 35428 566 35492
rect 582 35428 646 35492
rect 662 35428 726 35492
rect 422 35348 486 35412
rect 502 35348 566 35412
rect 582 35348 646 35412
rect 662 35348 726 35412
rect 422 35268 486 35332
rect 502 35268 566 35332
rect 582 35268 646 35332
rect 662 35268 726 35332
rect 422 35188 486 35252
rect 502 35188 566 35252
rect 582 35188 646 35252
rect 662 35188 726 35252
rect 2000 35428 2064 35492
rect 2080 35428 2144 35492
rect 2160 35428 2224 35492
rect 2240 35428 2304 35492
rect 2000 35348 2064 35412
rect 2080 35348 2144 35412
rect 2160 35348 2224 35412
rect 2240 35348 2304 35412
rect 2000 35268 2064 35332
rect 2080 35268 2144 35332
rect 2160 35268 2224 35332
rect 2240 35268 2304 35332
rect 2000 35188 2064 35252
rect 2080 35188 2144 35252
rect 2160 35188 2224 35252
rect 2240 35188 2304 35252
rect 50000 35428 50064 35492
rect 50080 35428 50144 35492
rect 50160 35428 50224 35492
rect 50240 35428 50304 35492
rect 50000 35348 50064 35412
rect 50080 35348 50144 35412
rect 50160 35348 50224 35412
rect 50240 35348 50304 35412
rect 50000 35268 50064 35332
rect 50080 35268 50144 35332
rect 50160 35268 50224 35332
rect 50240 35268 50304 35332
rect 50000 35188 50064 35252
rect 50080 35188 50144 35252
rect 50160 35188 50224 35252
rect 50240 35188 50304 35252
rect 62210 35428 62274 35492
rect 62290 35428 62354 35492
rect 62370 35428 62434 35492
rect 62450 35428 62514 35492
rect 62210 35348 62274 35412
rect 62290 35348 62354 35412
rect 62370 35348 62434 35412
rect 62450 35348 62514 35412
rect 62210 35268 62274 35332
rect 62290 35268 62354 35332
rect 62370 35268 62434 35332
rect 62450 35268 62514 35332
rect 65260 35388 65324 35392
rect 65260 35332 65264 35388
rect 65264 35332 65320 35388
rect 65320 35332 65324 35388
rect 65260 35328 65324 35332
rect 65340 35388 65404 35392
rect 65340 35332 65344 35388
rect 65344 35332 65400 35388
rect 65400 35332 65404 35388
rect 65340 35328 65404 35332
rect 65420 35388 65484 35392
rect 65420 35332 65424 35388
rect 65424 35332 65480 35388
rect 65480 35332 65484 35388
rect 65420 35328 65484 35332
rect 65500 35388 65564 35392
rect 65500 35332 65504 35388
rect 65504 35332 65560 35388
rect 65560 35332 65564 35388
rect 65500 35328 65564 35332
rect 62210 35188 62274 35252
rect 62290 35188 62354 35252
rect 62370 35188 62434 35252
rect 62450 35188 62514 35252
rect 63724 34988 63788 35052
rect 1118 34732 1182 34796
rect 1198 34732 1262 34796
rect 1278 34732 1342 34796
rect 1358 34732 1422 34796
rect 1118 34652 1182 34716
rect 1198 34652 1262 34716
rect 1278 34652 1342 34716
rect 1358 34652 1422 34716
rect 1118 34572 1182 34636
rect 1198 34572 1262 34636
rect 1278 34572 1342 34636
rect 1358 34572 1422 34636
rect 1118 34492 1182 34556
rect 1198 34492 1262 34556
rect 1278 34492 1342 34556
rect 1358 34492 1422 34556
rect 2920 34732 2984 34796
rect 3000 34732 3064 34796
rect 3080 34732 3144 34796
rect 3160 34732 3224 34796
rect 2920 34652 2984 34716
rect 3000 34652 3064 34716
rect 3080 34652 3144 34716
rect 3160 34652 3224 34716
rect 2920 34572 2984 34636
rect 3000 34572 3064 34636
rect 3080 34572 3144 34636
rect 3160 34572 3224 34636
rect 2920 34492 2984 34556
rect 3000 34492 3064 34556
rect 3080 34492 3144 34556
rect 3160 34492 3224 34556
rect 50920 34732 50984 34796
rect 51000 34732 51064 34796
rect 51080 34732 51144 34796
rect 51160 34732 51224 34796
rect 50920 34652 50984 34716
rect 51000 34652 51064 34716
rect 51080 34652 51144 34716
rect 51160 34652 51224 34716
rect 50920 34572 50984 34636
rect 51000 34572 51064 34636
rect 51080 34572 51144 34636
rect 51160 34572 51224 34636
rect 50920 34492 50984 34556
rect 51000 34492 51064 34556
rect 51080 34492 51144 34556
rect 51160 34492 51224 34556
rect 61514 34732 61578 34796
rect 61594 34732 61658 34796
rect 61674 34732 61738 34796
rect 61754 34732 61818 34796
rect 64340 34844 64404 34848
rect 64340 34788 64344 34844
rect 64344 34788 64400 34844
rect 64400 34788 64404 34844
rect 64340 34784 64404 34788
rect 64420 34844 64484 34848
rect 64420 34788 64424 34844
rect 64424 34788 64480 34844
rect 64480 34788 64484 34844
rect 64420 34784 64484 34788
rect 64500 34844 64564 34848
rect 64500 34788 64504 34844
rect 64504 34788 64560 34844
rect 64560 34788 64564 34844
rect 64500 34784 64564 34788
rect 64580 34844 64644 34848
rect 64580 34788 64584 34844
rect 64584 34788 64640 34844
rect 64640 34788 64644 34844
rect 64580 34784 64644 34788
rect 61514 34652 61578 34716
rect 61594 34652 61658 34716
rect 61674 34652 61738 34716
rect 61754 34652 61818 34716
rect 61514 34572 61578 34636
rect 61594 34572 61658 34636
rect 61674 34572 61738 34636
rect 61754 34572 61818 34636
rect 61514 34492 61578 34556
rect 61594 34492 61658 34556
rect 61674 34492 61738 34556
rect 61754 34492 61818 34556
rect 65260 34300 65324 34304
rect 65260 34244 65264 34300
rect 65264 34244 65320 34300
rect 65320 34244 65324 34300
rect 65260 34240 65324 34244
rect 65340 34300 65404 34304
rect 65340 34244 65344 34300
rect 65344 34244 65400 34300
rect 65400 34244 65404 34300
rect 65340 34240 65404 34244
rect 65420 34300 65484 34304
rect 65420 34244 65424 34300
rect 65424 34244 65480 34300
rect 65480 34244 65484 34300
rect 65420 34240 65484 34244
rect 65500 34300 65564 34304
rect 65500 34244 65504 34300
rect 65504 34244 65560 34300
rect 65560 34244 65564 34300
rect 65500 34240 65564 34244
rect 64340 33756 64404 33760
rect 64340 33700 64344 33756
rect 64344 33700 64400 33756
rect 64400 33700 64404 33756
rect 64340 33696 64404 33700
rect 64420 33756 64484 33760
rect 64420 33700 64424 33756
rect 64424 33700 64480 33756
rect 64480 33700 64484 33756
rect 64420 33696 64484 33700
rect 64500 33756 64564 33760
rect 64500 33700 64504 33756
rect 64504 33700 64560 33756
rect 64560 33700 64564 33756
rect 64500 33696 64564 33700
rect 64580 33756 64644 33760
rect 64580 33700 64584 33756
rect 64584 33700 64640 33756
rect 64640 33700 64644 33756
rect 64580 33696 64644 33700
rect 65260 33212 65324 33216
rect 65260 33156 65264 33212
rect 65264 33156 65320 33212
rect 65320 33156 65324 33212
rect 65260 33152 65324 33156
rect 65340 33212 65404 33216
rect 65340 33156 65344 33212
rect 65344 33156 65400 33212
rect 65400 33156 65404 33212
rect 65340 33152 65404 33156
rect 65420 33212 65484 33216
rect 65420 33156 65424 33212
rect 65424 33156 65480 33212
rect 65480 33156 65484 33212
rect 65420 33152 65484 33156
rect 65500 33212 65564 33216
rect 65500 33156 65504 33212
rect 65504 33156 65560 33212
rect 65560 33156 65564 33212
rect 65500 33152 65564 33156
rect 63908 33084 63972 33148
rect 64340 32668 64404 32672
rect 64340 32612 64344 32668
rect 64344 32612 64400 32668
rect 64400 32612 64404 32668
rect 64340 32608 64404 32612
rect 64420 32668 64484 32672
rect 64420 32612 64424 32668
rect 64424 32612 64480 32668
rect 64480 32612 64484 32668
rect 64420 32608 64484 32612
rect 64500 32668 64564 32672
rect 64500 32612 64504 32668
rect 64504 32612 64560 32668
rect 64560 32612 64564 32668
rect 64500 32608 64564 32612
rect 64580 32668 64644 32672
rect 64580 32612 64584 32668
rect 64584 32612 64640 32668
rect 64640 32612 64644 32668
rect 64580 32608 64644 32612
rect 64092 32404 64156 32468
rect 65260 32124 65324 32128
rect 65260 32068 65264 32124
rect 65264 32068 65320 32124
rect 65320 32068 65324 32124
rect 65260 32064 65324 32068
rect 65340 32124 65404 32128
rect 65340 32068 65344 32124
rect 65344 32068 65400 32124
rect 65400 32068 65404 32124
rect 65340 32064 65404 32068
rect 65420 32124 65484 32128
rect 65420 32068 65424 32124
rect 65424 32068 65480 32124
rect 65480 32068 65484 32124
rect 65420 32064 65484 32068
rect 65500 32124 65564 32128
rect 65500 32068 65504 32124
rect 65504 32068 65560 32124
rect 65560 32068 65564 32124
rect 65500 32064 65564 32068
rect 64340 31580 64404 31584
rect 64340 31524 64344 31580
rect 64344 31524 64400 31580
rect 64400 31524 64404 31580
rect 64340 31520 64404 31524
rect 64420 31580 64484 31584
rect 64420 31524 64424 31580
rect 64424 31524 64480 31580
rect 64480 31524 64484 31580
rect 64420 31520 64484 31524
rect 64500 31580 64564 31584
rect 64500 31524 64504 31580
rect 64504 31524 64560 31580
rect 64560 31524 64564 31580
rect 64500 31520 64564 31524
rect 64580 31580 64644 31584
rect 64580 31524 64584 31580
rect 64584 31524 64640 31580
rect 64640 31524 64644 31580
rect 64580 31520 64644 31524
rect 65260 31036 65324 31040
rect 65260 30980 65264 31036
rect 65264 30980 65320 31036
rect 65320 30980 65324 31036
rect 65260 30976 65324 30980
rect 65340 31036 65404 31040
rect 65340 30980 65344 31036
rect 65344 30980 65400 31036
rect 65400 30980 65404 31036
rect 65340 30976 65404 30980
rect 65420 31036 65484 31040
rect 65420 30980 65424 31036
rect 65424 30980 65480 31036
rect 65480 30980 65484 31036
rect 65420 30976 65484 30980
rect 65500 31036 65564 31040
rect 65500 30980 65504 31036
rect 65504 30980 65560 31036
rect 65560 30980 65564 31036
rect 65500 30976 65564 30980
rect 64340 30492 64404 30496
rect 64340 30436 64344 30492
rect 64344 30436 64400 30492
rect 64400 30436 64404 30492
rect 64340 30432 64404 30436
rect 64420 30492 64484 30496
rect 64420 30436 64424 30492
rect 64424 30436 64480 30492
rect 64480 30436 64484 30492
rect 64420 30432 64484 30436
rect 64500 30492 64564 30496
rect 64500 30436 64504 30492
rect 64504 30436 64560 30492
rect 64560 30436 64564 30492
rect 64500 30432 64564 30436
rect 64580 30492 64644 30496
rect 64580 30436 64584 30492
rect 64584 30436 64640 30492
rect 64640 30436 64644 30492
rect 64580 30432 64644 30436
rect 65260 29948 65324 29952
rect 65260 29892 65264 29948
rect 65264 29892 65320 29948
rect 65320 29892 65324 29948
rect 65260 29888 65324 29892
rect 65340 29948 65404 29952
rect 65340 29892 65344 29948
rect 65344 29892 65400 29948
rect 65400 29892 65404 29948
rect 65340 29888 65404 29892
rect 65420 29948 65484 29952
rect 65420 29892 65424 29948
rect 65424 29892 65480 29948
rect 65480 29892 65484 29948
rect 65420 29888 65484 29892
rect 65500 29948 65564 29952
rect 65500 29892 65504 29948
rect 65504 29892 65560 29948
rect 65560 29892 65564 29948
rect 65500 29888 65564 29892
rect 64340 29404 64404 29408
rect 64340 29348 64344 29404
rect 64344 29348 64400 29404
rect 64400 29348 64404 29404
rect 64340 29344 64404 29348
rect 64420 29404 64484 29408
rect 64420 29348 64424 29404
rect 64424 29348 64480 29404
rect 64480 29348 64484 29404
rect 64420 29344 64484 29348
rect 64500 29404 64564 29408
rect 64500 29348 64504 29404
rect 64504 29348 64560 29404
rect 64560 29348 64564 29404
rect 64500 29344 64564 29348
rect 64580 29404 64644 29408
rect 64580 29348 64584 29404
rect 64584 29348 64640 29404
rect 64640 29348 64644 29404
rect 64580 29344 64644 29348
rect 65260 28860 65324 28864
rect 65260 28804 65264 28860
rect 65264 28804 65320 28860
rect 65320 28804 65324 28860
rect 65260 28800 65324 28804
rect 65340 28860 65404 28864
rect 65340 28804 65344 28860
rect 65344 28804 65400 28860
rect 65400 28804 65404 28860
rect 65340 28800 65404 28804
rect 65420 28860 65484 28864
rect 65420 28804 65424 28860
rect 65424 28804 65480 28860
rect 65480 28804 65484 28860
rect 65420 28800 65484 28804
rect 65500 28860 65564 28864
rect 65500 28804 65504 28860
rect 65504 28804 65560 28860
rect 65560 28804 65564 28860
rect 65500 28800 65564 28804
rect 64340 28316 64404 28320
rect 64340 28260 64344 28316
rect 64344 28260 64400 28316
rect 64400 28260 64404 28316
rect 64340 28256 64404 28260
rect 64420 28316 64484 28320
rect 64420 28260 64424 28316
rect 64424 28260 64480 28316
rect 64480 28260 64484 28316
rect 64420 28256 64484 28260
rect 64500 28316 64564 28320
rect 64500 28260 64504 28316
rect 64504 28260 64560 28316
rect 64560 28260 64564 28316
rect 64500 28256 64564 28260
rect 64580 28316 64644 28320
rect 64580 28260 64584 28316
rect 64584 28260 64640 28316
rect 64640 28260 64644 28316
rect 64580 28256 64644 28260
rect 65260 27772 65324 27776
rect 65260 27716 65264 27772
rect 65264 27716 65320 27772
rect 65320 27716 65324 27772
rect 65260 27712 65324 27716
rect 65340 27772 65404 27776
rect 65340 27716 65344 27772
rect 65344 27716 65400 27772
rect 65400 27716 65404 27772
rect 65340 27712 65404 27716
rect 65420 27772 65484 27776
rect 65420 27716 65424 27772
rect 65424 27716 65480 27772
rect 65480 27716 65484 27772
rect 65420 27712 65484 27716
rect 65500 27772 65564 27776
rect 65500 27716 65504 27772
rect 65504 27716 65560 27772
rect 65560 27716 65564 27772
rect 65500 27712 65564 27716
rect 64340 27228 64404 27232
rect 64340 27172 64344 27228
rect 64344 27172 64400 27228
rect 64400 27172 64404 27228
rect 64340 27168 64404 27172
rect 64420 27228 64484 27232
rect 64420 27172 64424 27228
rect 64424 27172 64480 27228
rect 64480 27172 64484 27228
rect 64420 27168 64484 27172
rect 64500 27228 64564 27232
rect 64500 27172 64504 27228
rect 64504 27172 64560 27228
rect 64560 27172 64564 27228
rect 64500 27168 64564 27172
rect 64580 27228 64644 27232
rect 64580 27172 64584 27228
rect 64584 27172 64640 27228
rect 64640 27172 64644 27228
rect 64580 27168 64644 27172
rect 65260 26684 65324 26688
rect 65260 26628 65264 26684
rect 65264 26628 65320 26684
rect 65320 26628 65324 26684
rect 65260 26624 65324 26628
rect 65340 26684 65404 26688
rect 65340 26628 65344 26684
rect 65344 26628 65400 26684
rect 65400 26628 65404 26684
rect 65340 26624 65404 26628
rect 65420 26684 65484 26688
rect 65420 26628 65424 26684
rect 65424 26628 65480 26684
rect 65480 26628 65484 26684
rect 65420 26624 65484 26628
rect 65500 26684 65564 26688
rect 65500 26628 65504 26684
rect 65504 26628 65560 26684
rect 65560 26628 65564 26684
rect 65500 26624 65564 26628
rect 64340 26140 64404 26144
rect 64340 26084 64344 26140
rect 64344 26084 64400 26140
rect 64400 26084 64404 26140
rect 64340 26080 64404 26084
rect 64420 26140 64484 26144
rect 64420 26084 64424 26140
rect 64424 26084 64480 26140
rect 64480 26084 64484 26140
rect 64420 26080 64484 26084
rect 64500 26140 64564 26144
rect 64500 26084 64504 26140
rect 64504 26084 64560 26140
rect 64560 26084 64564 26140
rect 64500 26080 64564 26084
rect 64580 26140 64644 26144
rect 64580 26084 64584 26140
rect 64584 26084 64640 26140
rect 64640 26084 64644 26140
rect 64580 26080 64644 26084
rect 65260 25596 65324 25600
rect 65260 25540 65264 25596
rect 65264 25540 65320 25596
rect 65320 25540 65324 25596
rect 65260 25536 65324 25540
rect 65340 25596 65404 25600
rect 65340 25540 65344 25596
rect 65344 25540 65400 25596
rect 65400 25540 65404 25596
rect 65340 25536 65404 25540
rect 65420 25596 65484 25600
rect 65420 25540 65424 25596
rect 65424 25540 65480 25596
rect 65480 25540 65484 25596
rect 65420 25536 65484 25540
rect 65500 25596 65564 25600
rect 65500 25540 65504 25596
rect 65504 25540 65560 25596
rect 65560 25540 65564 25596
rect 65500 25536 65564 25540
rect 64340 25052 64404 25056
rect 64340 24996 64344 25052
rect 64344 24996 64400 25052
rect 64400 24996 64404 25052
rect 64340 24992 64404 24996
rect 64420 25052 64484 25056
rect 64420 24996 64424 25052
rect 64424 24996 64480 25052
rect 64480 24996 64484 25052
rect 64420 24992 64484 24996
rect 64500 25052 64564 25056
rect 64500 24996 64504 25052
rect 64504 24996 64560 25052
rect 64560 24996 64564 25052
rect 64500 24992 64564 24996
rect 64580 25052 64644 25056
rect 64580 24996 64584 25052
rect 64584 24996 64640 25052
rect 64640 24996 64644 25052
rect 64580 24992 64644 24996
rect 65260 24508 65324 24512
rect 65260 24452 65264 24508
rect 65264 24452 65320 24508
rect 65320 24452 65324 24508
rect 65260 24448 65324 24452
rect 65340 24508 65404 24512
rect 65340 24452 65344 24508
rect 65344 24452 65400 24508
rect 65400 24452 65404 24508
rect 65340 24448 65404 24452
rect 65420 24508 65484 24512
rect 65420 24452 65424 24508
rect 65424 24452 65480 24508
rect 65480 24452 65484 24508
rect 65420 24448 65484 24452
rect 65500 24508 65564 24512
rect 65500 24452 65504 24508
rect 65504 24452 65560 24508
rect 65560 24452 65564 24508
rect 65500 24448 65564 24452
rect 64340 23964 64404 23968
rect 64340 23908 64344 23964
rect 64344 23908 64400 23964
rect 64400 23908 64404 23964
rect 64340 23904 64404 23908
rect 64420 23964 64484 23968
rect 64420 23908 64424 23964
rect 64424 23908 64480 23964
rect 64480 23908 64484 23964
rect 64420 23904 64484 23908
rect 64500 23964 64564 23968
rect 64500 23908 64504 23964
rect 64504 23908 64560 23964
rect 64560 23908 64564 23964
rect 64500 23904 64564 23908
rect 64580 23964 64644 23968
rect 64580 23908 64584 23964
rect 64584 23908 64640 23964
rect 64640 23908 64644 23964
rect 64580 23904 64644 23908
rect 65260 23420 65324 23424
rect 65260 23364 65264 23420
rect 65264 23364 65320 23420
rect 65320 23364 65324 23420
rect 65260 23360 65324 23364
rect 65340 23420 65404 23424
rect 65340 23364 65344 23420
rect 65344 23364 65400 23420
rect 65400 23364 65404 23420
rect 65340 23360 65404 23364
rect 65420 23420 65484 23424
rect 65420 23364 65424 23420
rect 65424 23364 65480 23420
rect 65480 23364 65484 23420
rect 65420 23360 65484 23364
rect 65500 23420 65564 23424
rect 65500 23364 65504 23420
rect 65504 23364 65560 23420
rect 65560 23364 65564 23420
rect 65500 23360 65564 23364
rect 64340 22876 64404 22880
rect 64340 22820 64344 22876
rect 64344 22820 64400 22876
rect 64400 22820 64404 22876
rect 64340 22816 64404 22820
rect 64420 22876 64484 22880
rect 64420 22820 64424 22876
rect 64424 22820 64480 22876
rect 64480 22820 64484 22876
rect 64420 22816 64484 22820
rect 64500 22876 64564 22880
rect 64500 22820 64504 22876
rect 64504 22820 64560 22876
rect 64560 22820 64564 22876
rect 64500 22816 64564 22820
rect 64580 22876 64644 22880
rect 64580 22820 64584 22876
rect 64584 22820 64640 22876
rect 64640 22820 64644 22876
rect 64580 22816 64644 22820
rect 65260 22332 65324 22336
rect 65260 22276 65264 22332
rect 65264 22276 65320 22332
rect 65320 22276 65324 22332
rect 65260 22272 65324 22276
rect 65340 22332 65404 22336
rect 65340 22276 65344 22332
rect 65344 22276 65400 22332
rect 65400 22276 65404 22332
rect 65340 22272 65404 22276
rect 65420 22332 65484 22336
rect 65420 22276 65424 22332
rect 65424 22276 65480 22332
rect 65480 22276 65484 22332
rect 65420 22272 65484 22276
rect 65500 22332 65564 22336
rect 65500 22276 65504 22332
rect 65504 22276 65560 22332
rect 65560 22276 65564 22332
rect 65500 22272 65564 22276
rect 64340 21788 64404 21792
rect 64340 21732 64344 21788
rect 64344 21732 64400 21788
rect 64400 21732 64404 21788
rect 64340 21728 64404 21732
rect 64420 21788 64484 21792
rect 64420 21732 64424 21788
rect 64424 21732 64480 21788
rect 64480 21732 64484 21788
rect 64420 21728 64484 21732
rect 64500 21788 64564 21792
rect 64500 21732 64504 21788
rect 64504 21732 64560 21788
rect 64560 21732 64564 21788
rect 64500 21728 64564 21732
rect 64580 21788 64644 21792
rect 64580 21732 64584 21788
rect 64584 21732 64640 21788
rect 64640 21732 64644 21788
rect 64580 21728 64644 21732
rect 65260 21244 65324 21248
rect 65260 21188 65264 21244
rect 65264 21188 65320 21244
rect 65320 21188 65324 21244
rect 65260 21184 65324 21188
rect 65340 21244 65404 21248
rect 65340 21188 65344 21244
rect 65344 21188 65400 21244
rect 65400 21188 65404 21244
rect 65340 21184 65404 21188
rect 65420 21244 65484 21248
rect 65420 21188 65424 21244
rect 65424 21188 65480 21244
rect 65480 21188 65484 21244
rect 65420 21184 65484 21188
rect 65500 21244 65564 21248
rect 65500 21188 65504 21244
rect 65504 21188 65560 21244
rect 65560 21188 65564 21244
rect 65500 21184 65564 21188
rect 64340 20700 64404 20704
rect 64340 20644 64344 20700
rect 64344 20644 64400 20700
rect 64400 20644 64404 20700
rect 64340 20640 64404 20644
rect 64420 20700 64484 20704
rect 64420 20644 64424 20700
rect 64424 20644 64480 20700
rect 64480 20644 64484 20700
rect 64420 20640 64484 20644
rect 64500 20700 64564 20704
rect 64500 20644 64504 20700
rect 64504 20644 64560 20700
rect 64560 20644 64564 20700
rect 64500 20640 64564 20644
rect 64580 20700 64644 20704
rect 64580 20644 64584 20700
rect 64584 20644 64640 20700
rect 64640 20644 64644 20700
rect 64580 20640 64644 20644
rect 65260 20156 65324 20160
rect 65260 20100 65264 20156
rect 65264 20100 65320 20156
rect 65320 20100 65324 20156
rect 65260 20096 65324 20100
rect 65340 20156 65404 20160
rect 65340 20100 65344 20156
rect 65344 20100 65400 20156
rect 65400 20100 65404 20156
rect 65340 20096 65404 20100
rect 65420 20156 65484 20160
rect 65420 20100 65424 20156
rect 65424 20100 65480 20156
rect 65480 20100 65484 20156
rect 65420 20096 65484 20100
rect 65500 20156 65564 20160
rect 65500 20100 65504 20156
rect 65504 20100 65560 20156
rect 65560 20100 65564 20156
rect 65500 20096 65564 20100
rect 64340 19612 64404 19616
rect 64340 19556 64344 19612
rect 64344 19556 64400 19612
rect 64400 19556 64404 19612
rect 64340 19552 64404 19556
rect 64420 19612 64484 19616
rect 64420 19556 64424 19612
rect 64424 19556 64480 19612
rect 64480 19556 64484 19612
rect 64420 19552 64484 19556
rect 64500 19612 64564 19616
rect 64500 19556 64504 19612
rect 64504 19556 64560 19612
rect 64560 19556 64564 19612
rect 64500 19552 64564 19556
rect 64580 19612 64644 19616
rect 64580 19556 64584 19612
rect 64584 19556 64640 19612
rect 64640 19556 64644 19612
rect 64580 19552 64644 19556
rect 65260 19068 65324 19072
rect 65260 19012 65264 19068
rect 65264 19012 65320 19068
rect 65320 19012 65324 19068
rect 65260 19008 65324 19012
rect 65340 19068 65404 19072
rect 65340 19012 65344 19068
rect 65344 19012 65400 19068
rect 65400 19012 65404 19068
rect 65340 19008 65404 19012
rect 65420 19068 65484 19072
rect 65420 19012 65424 19068
rect 65424 19012 65480 19068
rect 65480 19012 65484 19068
rect 65420 19008 65484 19012
rect 65500 19068 65564 19072
rect 65500 19012 65504 19068
rect 65504 19012 65560 19068
rect 65560 19012 65564 19068
rect 65500 19008 65564 19012
rect 64340 18524 64404 18528
rect 64340 18468 64344 18524
rect 64344 18468 64400 18524
rect 64400 18468 64404 18524
rect 64340 18464 64404 18468
rect 64420 18524 64484 18528
rect 64420 18468 64424 18524
rect 64424 18468 64480 18524
rect 64480 18468 64484 18524
rect 64420 18464 64484 18468
rect 64500 18524 64564 18528
rect 64500 18468 64504 18524
rect 64504 18468 64560 18524
rect 64560 18468 64564 18524
rect 64500 18464 64564 18468
rect 64580 18524 64644 18528
rect 64580 18468 64584 18524
rect 64584 18468 64640 18524
rect 64640 18468 64644 18524
rect 64580 18464 64644 18468
rect 65260 17980 65324 17984
rect 65260 17924 65264 17980
rect 65264 17924 65320 17980
rect 65320 17924 65324 17980
rect 65260 17920 65324 17924
rect 65340 17980 65404 17984
rect 65340 17924 65344 17980
rect 65344 17924 65400 17980
rect 65400 17924 65404 17980
rect 65340 17920 65404 17924
rect 65420 17980 65484 17984
rect 65420 17924 65424 17980
rect 65424 17924 65480 17980
rect 65480 17924 65484 17980
rect 65420 17920 65484 17924
rect 65500 17980 65564 17984
rect 65500 17924 65504 17980
rect 65504 17924 65560 17980
rect 65560 17924 65564 17980
rect 65500 17920 65564 17924
rect 63724 17852 63788 17916
rect 64340 17436 64404 17440
rect 64340 17380 64344 17436
rect 64344 17380 64400 17436
rect 64400 17380 64404 17436
rect 64340 17376 64404 17380
rect 64420 17436 64484 17440
rect 64420 17380 64424 17436
rect 64424 17380 64480 17436
rect 64480 17380 64484 17436
rect 64420 17376 64484 17380
rect 64500 17436 64564 17440
rect 64500 17380 64504 17436
rect 64504 17380 64560 17436
rect 64560 17380 64564 17436
rect 64500 17376 64564 17380
rect 64580 17436 64644 17440
rect 64580 17380 64584 17436
rect 64584 17380 64640 17436
rect 64640 17380 64644 17436
rect 64580 17376 64644 17380
rect 62804 17172 62868 17236
rect 65260 16892 65324 16896
rect 65260 16836 65264 16892
rect 65264 16836 65320 16892
rect 65320 16836 65324 16892
rect 65260 16832 65324 16836
rect 65340 16892 65404 16896
rect 65340 16836 65344 16892
rect 65344 16836 65400 16892
rect 65400 16836 65404 16892
rect 65340 16832 65404 16836
rect 65420 16892 65484 16896
rect 65420 16836 65424 16892
rect 65424 16836 65480 16892
rect 65480 16836 65484 16892
rect 65420 16832 65484 16836
rect 65500 16892 65564 16896
rect 65500 16836 65504 16892
rect 65504 16836 65560 16892
rect 65560 16836 65564 16892
rect 65500 16832 65564 16836
rect 64340 16348 64404 16352
rect 64340 16292 64344 16348
rect 64344 16292 64400 16348
rect 64400 16292 64404 16348
rect 64340 16288 64404 16292
rect 64420 16348 64484 16352
rect 64420 16292 64424 16348
rect 64424 16292 64480 16348
rect 64480 16292 64484 16348
rect 64420 16288 64484 16292
rect 64500 16348 64564 16352
rect 64500 16292 64504 16348
rect 64504 16292 64560 16348
rect 64560 16292 64564 16348
rect 64500 16288 64564 16292
rect 64580 16348 64644 16352
rect 64580 16292 64584 16348
rect 64584 16292 64640 16348
rect 64640 16292 64644 16348
rect 64580 16288 64644 16292
rect 65260 15804 65324 15808
rect 65260 15748 65264 15804
rect 65264 15748 65320 15804
rect 65320 15748 65324 15804
rect 65260 15744 65324 15748
rect 65340 15804 65404 15808
rect 65340 15748 65344 15804
rect 65344 15748 65400 15804
rect 65400 15748 65404 15804
rect 65340 15744 65404 15748
rect 65420 15804 65484 15808
rect 65420 15748 65424 15804
rect 65424 15748 65480 15804
rect 65480 15748 65484 15804
rect 65420 15744 65484 15748
rect 65500 15804 65564 15808
rect 65500 15748 65504 15804
rect 65504 15748 65560 15804
rect 65560 15748 65564 15804
rect 65500 15744 65564 15748
rect 62620 15676 62684 15740
rect 64340 15260 64404 15264
rect 64340 15204 64344 15260
rect 64344 15204 64400 15260
rect 64400 15204 64404 15260
rect 64340 15200 64404 15204
rect 64420 15260 64484 15264
rect 64420 15204 64424 15260
rect 64424 15204 64480 15260
rect 64480 15204 64484 15260
rect 64420 15200 64484 15204
rect 64500 15260 64564 15264
rect 64500 15204 64504 15260
rect 64504 15204 64560 15260
rect 64560 15204 64564 15260
rect 64500 15200 64564 15204
rect 64580 15260 64644 15264
rect 64580 15204 64584 15260
rect 64584 15204 64640 15260
rect 64640 15204 64644 15260
rect 64580 15200 64644 15204
rect 65260 14716 65324 14720
rect 65260 14660 65264 14716
rect 65264 14660 65320 14716
rect 65320 14660 65324 14716
rect 65260 14656 65324 14660
rect 65340 14716 65404 14720
rect 65340 14660 65344 14716
rect 65344 14660 65400 14716
rect 65400 14660 65404 14716
rect 65340 14656 65404 14660
rect 65420 14716 65484 14720
rect 65420 14660 65424 14716
rect 65424 14660 65480 14716
rect 65480 14660 65484 14716
rect 65420 14656 65484 14660
rect 65500 14716 65564 14720
rect 65500 14660 65504 14716
rect 65504 14660 65560 14716
rect 65560 14660 65564 14716
rect 65500 14656 65564 14660
rect 64340 14172 64404 14176
rect 64340 14116 64344 14172
rect 64344 14116 64400 14172
rect 64400 14116 64404 14172
rect 64340 14112 64404 14116
rect 64420 14172 64484 14176
rect 64420 14116 64424 14172
rect 64424 14116 64480 14172
rect 64480 14116 64484 14172
rect 64420 14112 64484 14116
rect 64500 14172 64564 14176
rect 64500 14116 64504 14172
rect 64504 14116 64560 14172
rect 64560 14116 64564 14172
rect 64500 14112 64564 14116
rect 64580 14172 64644 14176
rect 64580 14116 64584 14172
rect 64584 14116 64640 14172
rect 64640 14116 64644 14172
rect 64580 14112 64644 14116
rect 65260 13628 65324 13632
rect 65260 13572 65264 13628
rect 65264 13572 65320 13628
rect 65320 13572 65324 13628
rect 65260 13568 65324 13572
rect 65340 13628 65404 13632
rect 65340 13572 65344 13628
rect 65344 13572 65400 13628
rect 65400 13572 65404 13628
rect 65340 13568 65404 13572
rect 65420 13628 65484 13632
rect 65420 13572 65424 13628
rect 65424 13572 65480 13628
rect 65480 13572 65484 13628
rect 65420 13568 65484 13572
rect 65500 13628 65564 13632
rect 65500 13572 65504 13628
rect 65504 13572 65560 13628
rect 65560 13572 65564 13628
rect 65500 13568 65564 13572
rect 64340 13084 64404 13088
rect 64340 13028 64344 13084
rect 64344 13028 64400 13084
rect 64400 13028 64404 13084
rect 64340 13024 64404 13028
rect 64420 13084 64484 13088
rect 64420 13028 64424 13084
rect 64424 13028 64480 13084
rect 64480 13028 64484 13084
rect 64420 13024 64484 13028
rect 64500 13084 64564 13088
rect 64500 13028 64504 13084
rect 64504 13028 64560 13084
rect 64560 13028 64564 13084
rect 64500 13024 64564 13028
rect 64580 13084 64644 13088
rect 64580 13028 64584 13084
rect 64584 13028 64640 13084
rect 64640 13028 64644 13084
rect 64580 13024 64644 13028
rect 65260 12540 65324 12544
rect 65260 12484 65264 12540
rect 65264 12484 65320 12540
rect 65320 12484 65324 12540
rect 65260 12480 65324 12484
rect 65340 12540 65404 12544
rect 65340 12484 65344 12540
rect 65344 12484 65400 12540
rect 65400 12484 65404 12540
rect 65340 12480 65404 12484
rect 65420 12540 65484 12544
rect 65420 12484 65424 12540
rect 65424 12484 65480 12540
rect 65480 12484 65484 12540
rect 65420 12480 65484 12484
rect 65500 12540 65564 12544
rect 65500 12484 65504 12540
rect 65504 12484 65560 12540
rect 65560 12484 65564 12540
rect 65500 12480 65564 12484
rect 64340 11996 64404 12000
rect 64340 11940 64344 11996
rect 64344 11940 64400 11996
rect 64400 11940 64404 11996
rect 64340 11936 64404 11940
rect 64420 11996 64484 12000
rect 64420 11940 64424 11996
rect 64424 11940 64480 11996
rect 64480 11940 64484 11996
rect 64420 11936 64484 11940
rect 64500 11996 64564 12000
rect 64500 11940 64504 11996
rect 64504 11940 64560 11996
rect 64560 11940 64564 11996
rect 64500 11936 64564 11940
rect 64580 11996 64644 12000
rect 64580 11940 64584 11996
rect 64584 11940 64640 11996
rect 64640 11940 64644 11996
rect 64580 11936 64644 11940
rect 65260 11452 65324 11456
rect 65260 11396 65264 11452
rect 65264 11396 65320 11452
rect 65320 11396 65324 11452
rect 65260 11392 65324 11396
rect 65340 11452 65404 11456
rect 65340 11396 65344 11452
rect 65344 11396 65400 11452
rect 65400 11396 65404 11452
rect 65340 11392 65404 11396
rect 65420 11452 65484 11456
rect 65420 11396 65424 11452
rect 65424 11396 65480 11452
rect 65480 11396 65484 11452
rect 65420 11392 65484 11396
rect 65500 11452 65564 11456
rect 65500 11396 65504 11452
rect 65504 11396 65560 11452
rect 65560 11396 65564 11452
rect 65500 11392 65564 11396
rect 64340 10908 64404 10912
rect 64340 10852 64344 10908
rect 64344 10852 64400 10908
rect 64400 10852 64404 10908
rect 64340 10848 64404 10852
rect 64420 10908 64484 10912
rect 64420 10852 64424 10908
rect 64424 10852 64480 10908
rect 64480 10852 64484 10908
rect 64420 10848 64484 10852
rect 64500 10908 64564 10912
rect 64500 10852 64504 10908
rect 64504 10852 64560 10908
rect 64560 10852 64564 10908
rect 64500 10848 64564 10852
rect 64580 10908 64644 10912
rect 64580 10852 64584 10908
rect 64584 10852 64640 10908
rect 64640 10852 64644 10908
rect 64580 10848 64644 10852
rect 65260 10364 65324 10368
rect 65260 10308 65264 10364
rect 65264 10308 65320 10364
rect 65320 10308 65324 10364
rect 65260 10304 65324 10308
rect 65340 10364 65404 10368
rect 65340 10308 65344 10364
rect 65344 10308 65400 10364
rect 65400 10308 65404 10364
rect 65340 10304 65404 10308
rect 65420 10364 65484 10368
rect 65420 10308 65424 10364
rect 65424 10308 65480 10364
rect 65480 10308 65484 10364
rect 65420 10304 65484 10308
rect 65500 10364 65564 10368
rect 65500 10308 65504 10364
rect 65504 10308 65560 10364
rect 65560 10308 65564 10364
rect 65500 10304 65564 10308
rect 64340 9820 64404 9824
rect 64340 9764 64344 9820
rect 64344 9764 64400 9820
rect 64400 9764 64404 9820
rect 64340 9760 64404 9764
rect 64420 9820 64484 9824
rect 64420 9764 64424 9820
rect 64424 9764 64480 9820
rect 64480 9764 64484 9820
rect 64420 9760 64484 9764
rect 64500 9820 64564 9824
rect 64500 9764 64504 9820
rect 64504 9764 64560 9820
rect 64560 9764 64564 9820
rect 64500 9760 64564 9764
rect 64580 9820 64644 9824
rect 64580 9764 64584 9820
rect 64584 9764 64640 9820
rect 64640 9764 64644 9820
rect 64580 9760 64644 9764
rect 65260 9276 65324 9280
rect 65260 9220 65264 9276
rect 65264 9220 65320 9276
rect 65320 9220 65324 9276
rect 65260 9216 65324 9220
rect 65340 9276 65404 9280
rect 65340 9220 65344 9276
rect 65344 9220 65400 9276
rect 65400 9220 65404 9276
rect 65340 9216 65404 9220
rect 65420 9276 65484 9280
rect 65420 9220 65424 9276
rect 65424 9220 65480 9276
rect 65480 9220 65484 9276
rect 65420 9216 65484 9220
rect 65500 9276 65564 9280
rect 65500 9220 65504 9276
rect 65504 9220 65560 9276
rect 65560 9220 65564 9276
rect 65500 9216 65564 9220
rect 64340 8732 64404 8736
rect 64340 8676 64344 8732
rect 64344 8676 64400 8732
rect 64400 8676 64404 8732
rect 64340 8672 64404 8676
rect 64420 8732 64484 8736
rect 64420 8676 64424 8732
rect 64424 8676 64480 8732
rect 64480 8676 64484 8732
rect 64420 8672 64484 8676
rect 64500 8732 64564 8736
rect 64500 8676 64504 8732
rect 64504 8676 64560 8732
rect 64560 8676 64564 8732
rect 64500 8672 64564 8676
rect 64580 8732 64644 8736
rect 64580 8676 64584 8732
rect 64584 8676 64640 8732
rect 64640 8676 64644 8732
rect 64580 8672 64644 8676
rect 65260 8188 65324 8192
rect 65260 8132 65264 8188
rect 65264 8132 65320 8188
rect 65320 8132 65324 8188
rect 65260 8128 65324 8132
rect 65340 8188 65404 8192
rect 65340 8132 65344 8188
rect 65344 8132 65400 8188
rect 65400 8132 65404 8188
rect 65340 8128 65404 8132
rect 65420 8188 65484 8192
rect 65420 8132 65424 8188
rect 65424 8132 65480 8188
rect 65480 8132 65484 8188
rect 65420 8128 65484 8132
rect 65500 8188 65564 8192
rect 65500 8132 65504 8188
rect 65504 8132 65560 8188
rect 65560 8132 65564 8188
rect 65500 8128 65564 8132
rect 64340 7644 64404 7648
rect 64340 7588 64344 7644
rect 64344 7588 64400 7644
rect 64400 7588 64404 7644
rect 64340 7584 64404 7588
rect 64420 7644 64484 7648
rect 64420 7588 64424 7644
rect 64424 7588 64480 7644
rect 64480 7588 64484 7644
rect 64420 7584 64484 7588
rect 64500 7644 64564 7648
rect 64500 7588 64504 7644
rect 64504 7588 64560 7644
rect 64560 7588 64564 7644
rect 64500 7584 64564 7588
rect 64580 7644 64644 7648
rect 64580 7588 64584 7644
rect 64584 7588 64640 7644
rect 64640 7588 64644 7644
rect 64580 7584 64644 7588
rect 63540 7380 63604 7444
rect 65260 7100 65324 7104
rect 65260 7044 65264 7100
rect 65264 7044 65320 7100
rect 65320 7044 65324 7100
rect 65260 7040 65324 7044
rect 65340 7100 65404 7104
rect 65340 7044 65344 7100
rect 65344 7044 65400 7100
rect 65400 7044 65404 7100
rect 65340 7040 65404 7044
rect 65420 7100 65484 7104
rect 65420 7044 65424 7100
rect 65424 7044 65480 7100
rect 65480 7044 65484 7100
rect 65420 7040 65484 7044
rect 65500 7100 65564 7104
rect 65500 7044 65504 7100
rect 65504 7044 65560 7100
rect 65560 7044 65564 7100
rect 65500 7040 65564 7044
rect 63908 6836 63972 6900
rect 64340 6556 64404 6560
rect 64340 6500 64344 6556
rect 64344 6500 64400 6556
rect 64400 6500 64404 6556
rect 64340 6496 64404 6500
rect 64420 6556 64484 6560
rect 64420 6500 64424 6556
rect 64424 6500 64480 6556
rect 64480 6500 64484 6556
rect 64420 6496 64484 6500
rect 64500 6556 64564 6560
rect 64500 6500 64504 6556
rect 64504 6500 64560 6556
rect 64560 6500 64564 6556
rect 64500 6496 64564 6500
rect 64580 6556 64644 6560
rect 64580 6500 64584 6556
rect 64584 6500 64640 6556
rect 64640 6500 64644 6556
rect 64580 6496 64644 6500
rect 65260 6012 65324 6016
rect 65260 5956 65264 6012
rect 65264 5956 65320 6012
rect 65320 5956 65324 6012
rect 65260 5952 65324 5956
rect 65340 6012 65404 6016
rect 65340 5956 65344 6012
rect 65344 5956 65400 6012
rect 65400 5956 65404 6012
rect 65340 5952 65404 5956
rect 65420 6012 65484 6016
rect 65420 5956 65424 6012
rect 65424 5956 65480 6012
rect 65480 5956 65484 6012
rect 65420 5952 65484 5956
rect 65500 6012 65564 6016
rect 65500 5956 65504 6012
rect 65504 5956 65560 6012
rect 65560 5956 65564 6012
rect 65500 5952 65564 5956
rect 64340 5468 64404 5472
rect 64340 5412 64344 5468
rect 64344 5412 64400 5468
rect 64400 5412 64404 5468
rect 64340 5408 64404 5412
rect 64420 5468 64484 5472
rect 64420 5412 64424 5468
rect 64424 5412 64480 5468
rect 64480 5412 64484 5468
rect 64420 5408 64484 5412
rect 64500 5468 64564 5472
rect 64500 5412 64504 5468
rect 64504 5412 64560 5468
rect 64560 5412 64564 5468
rect 64500 5408 64564 5412
rect 64580 5468 64644 5472
rect 64580 5412 64584 5468
rect 64584 5412 64640 5468
rect 64640 5412 64644 5468
rect 64580 5408 64644 5412
rect 65260 4924 65324 4928
rect 65260 4868 65264 4924
rect 65264 4868 65320 4924
rect 65320 4868 65324 4924
rect 65260 4864 65324 4868
rect 65340 4924 65404 4928
rect 65340 4868 65344 4924
rect 65344 4868 65400 4924
rect 65400 4868 65404 4924
rect 65340 4864 65404 4868
rect 65420 4924 65484 4928
rect 65420 4868 65424 4924
rect 65424 4868 65480 4924
rect 65480 4868 65484 4924
rect 65420 4864 65484 4868
rect 65500 4924 65564 4928
rect 65500 4868 65504 4924
rect 65504 4868 65560 4924
rect 65560 4868 65564 4924
rect 65500 4864 65564 4868
rect 64340 4380 64404 4384
rect 64340 4324 64344 4380
rect 64344 4324 64400 4380
rect 64400 4324 64404 4380
rect 64340 4320 64404 4324
rect 64420 4380 64484 4384
rect 64420 4324 64424 4380
rect 64424 4324 64480 4380
rect 64480 4324 64484 4380
rect 64420 4320 64484 4324
rect 64500 4380 64564 4384
rect 64500 4324 64504 4380
rect 64504 4324 64560 4380
rect 64560 4324 64564 4380
rect 64500 4320 64564 4324
rect 64580 4380 64644 4384
rect 64580 4324 64584 4380
rect 64584 4324 64640 4380
rect 64640 4324 64644 4380
rect 64580 4320 64644 4324
rect 65260 3836 65324 3840
rect 65260 3780 65264 3836
rect 65264 3780 65320 3836
rect 65320 3780 65324 3836
rect 65260 3776 65324 3780
rect 65340 3836 65404 3840
rect 65340 3780 65344 3836
rect 65344 3780 65400 3836
rect 65400 3780 65404 3836
rect 65340 3776 65404 3780
rect 65420 3836 65484 3840
rect 65420 3780 65424 3836
rect 65424 3780 65480 3836
rect 65480 3780 65484 3836
rect 65420 3776 65484 3780
rect 65500 3836 65564 3840
rect 65500 3780 65504 3836
rect 65504 3780 65560 3836
rect 65560 3780 65564 3836
rect 65500 3776 65564 3780
rect 64340 3292 64404 3296
rect 64340 3236 64344 3292
rect 64344 3236 64400 3292
rect 64400 3236 64404 3292
rect 64340 3232 64404 3236
rect 64420 3292 64484 3296
rect 64420 3236 64424 3292
rect 64424 3236 64480 3292
rect 64480 3236 64484 3292
rect 64420 3232 64484 3236
rect 64500 3292 64564 3296
rect 64500 3236 64504 3292
rect 64504 3236 64560 3292
rect 64560 3236 64564 3292
rect 64500 3232 64564 3236
rect 64580 3292 64644 3296
rect 64580 3236 64584 3292
rect 64584 3236 64640 3292
rect 64640 3236 64644 3292
rect 64580 3232 64644 3236
rect 1118 2958 1182 3022
rect 1198 2958 1262 3022
rect 1278 2958 1342 3022
rect 1358 2958 1422 3022
rect 1118 2878 1182 2942
rect 1198 2878 1262 2942
rect 1278 2878 1342 2942
rect 1358 2878 1422 2942
rect 1118 2798 1182 2862
rect 1198 2798 1262 2862
rect 1278 2798 1342 2862
rect 1358 2798 1422 2862
rect 1118 2718 1182 2782
rect 1198 2718 1262 2782
rect 1278 2718 1342 2782
rect 1358 2718 1422 2782
rect 61514 2958 61578 3022
rect 61594 2958 61658 3022
rect 61674 2958 61738 3022
rect 61754 2958 61818 3022
rect 61514 2878 61578 2942
rect 61594 2878 61658 2942
rect 61674 2878 61738 2942
rect 61754 2878 61818 2942
rect 61514 2798 61578 2862
rect 61594 2798 61658 2862
rect 61674 2798 61738 2862
rect 61754 2798 61818 2862
rect 61514 2718 61578 2782
rect 61594 2718 61658 2782
rect 61674 2718 61738 2782
rect 61754 2718 61818 2782
rect 65260 2748 65324 2752
rect 65260 2692 65264 2748
rect 65264 2692 65320 2748
rect 65320 2692 65324 2748
rect 65260 2688 65324 2692
rect 65340 2748 65404 2752
rect 65340 2692 65344 2748
rect 65344 2692 65400 2748
rect 65400 2692 65404 2748
rect 65340 2688 65404 2692
rect 65420 2748 65484 2752
rect 65420 2692 65424 2748
rect 65424 2692 65480 2748
rect 65480 2692 65484 2748
rect 65420 2688 65484 2692
rect 65500 2748 65564 2752
rect 65500 2692 65504 2748
rect 65504 2692 65560 2748
rect 65560 2692 65564 2748
rect 65500 2688 65564 2692
rect 422 2262 486 2326
rect 502 2262 566 2326
rect 582 2262 646 2326
rect 662 2262 726 2326
rect 422 2182 486 2246
rect 502 2182 566 2246
rect 582 2182 646 2246
rect 662 2182 726 2246
rect 422 2102 486 2166
rect 502 2102 566 2166
rect 582 2102 646 2166
rect 662 2102 726 2166
rect 422 2022 486 2086
rect 502 2022 566 2086
rect 582 2022 646 2086
rect 662 2022 726 2086
rect 62210 2262 62274 2326
rect 62290 2262 62354 2326
rect 62370 2262 62434 2326
rect 62450 2262 62514 2326
rect 62210 2182 62274 2246
rect 62290 2182 62354 2246
rect 62370 2182 62434 2246
rect 62450 2182 62514 2246
rect 62210 2102 62274 2166
rect 62290 2102 62354 2166
rect 62370 2102 62434 2166
rect 62450 2102 62514 2166
rect 64340 2204 64404 2208
rect 64340 2148 64344 2204
rect 64344 2148 64400 2204
rect 64400 2148 64404 2204
rect 64340 2144 64404 2148
rect 64420 2204 64484 2208
rect 64420 2148 64424 2204
rect 64424 2148 64480 2204
rect 64480 2148 64484 2204
rect 64420 2144 64484 2148
rect 64500 2204 64564 2208
rect 64500 2148 64504 2204
rect 64504 2148 64560 2204
rect 64560 2148 64564 2204
rect 64500 2144 64564 2148
rect 64580 2204 64644 2208
rect 64580 2148 64584 2204
rect 64584 2148 64640 2204
rect 64640 2148 64644 2204
rect 64580 2144 64644 2148
rect 62210 2022 62274 2086
rect 62290 2022 62354 2086
rect 62370 2022 62434 2086
rect 62450 2022 62514 2086
rect 48941 1864 49005 1868
rect 48941 1808 48962 1864
rect 48962 1808 49005 1864
rect 48941 1804 49005 1808
rect 49372 1804 49436 1868
rect 49674 1728 49738 1732
rect 49674 1672 49698 1728
rect 49698 1672 49738 1728
rect 49674 1668 49738 1672
rect 49079 1532 49143 1596
rect 49217 1532 49281 1596
rect 65260 1660 65324 1664
rect 65260 1604 65264 1660
rect 65264 1604 65320 1660
rect 65320 1604 65324 1660
rect 65260 1600 65324 1604
rect 65340 1660 65404 1664
rect 65340 1604 65344 1660
rect 65344 1604 65400 1660
rect 65400 1604 65404 1660
rect 65340 1600 65404 1604
rect 65420 1660 65484 1664
rect 65420 1604 65424 1660
rect 65424 1604 65480 1660
rect 65480 1604 65484 1660
rect 65420 1600 65484 1604
rect 65500 1660 65564 1664
rect 65500 1604 65504 1660
rect 65504 1604 65560 1660
rect 65560 1604 65564 1660
rect 65500 1600 65564 1604
rect 49924 1260 49988 1324
rect 64340 1116 64404 1120
rect 64340 1060 64344 1116
rect 64344 1060 64400 1116
rect 64400 1060 64404 1116
rect 64340 1056 64404 1060
rect 64420 1116 64484 1120
rect 64420 1060 64424 1116
rect 64424 1060 64480 1116
rect 64480 1060 64484 1116
rect 64420 1056 64484 1060
rect 64500 1116 64564 1120
rect 64500 1060 64504 1116
rect 64504 1060 64560 1116
rect 64560 1060 64564 1116
rect 64500 1056 64564 1060
rect 64580 1116 64644 1120
rect 64580 1060 64584 1116
rect 64584 1060 64640 1116
rect 64640 1060 64644 1116
rect 64580 1056 64644 1060
rect 65260 572 65324 576
rect 65260 516 65264 572
rect 65264 516 65320 572
rect 65320 516 65324 572
rect 65260 512 65324 516
rect 65340 572 65404 576
rect 65340 516 65344 572
rect 65344 516 65400 572
rect 65400 516 65404 572
rect 65340 512 65404 516
rect 65420 572 65484 576
rect 65420 516 65424 572
rect 65424 516 65480 572
rect 65480 516 65484 572
rect 65420 512 65484 516
rect 65500 572 65564 576
rect 65500 516 65504 572
rect 65504 516 65560 572
rect 65560 516 65564 572
rect 65500 512 65564 516
<< metal4 >>
rect 1992 44640 2312 44656
rect 1992 44576 2000 44640
rect 2064 44576 2080 44640
rect 2144 44576 2160 44640
rect 2224 44576 2240 44640
rect 2304 44576 2312 44640
rect 1992 43552 2312 44576
rect 1992 43488 2000 43552
rect 2064 43488 2080 43552
rect 2144 43488 2160 43552
rect 2224 43488 2240 43552
rect 2304 43488 2312 43552
rect 1992 42464 2312 43488
rect 1992 42400 2000 42464
rect 2064 42400 2080 42464
rect 2144 42400 2160 42464
rect 2224 42400 2240 42464
rect 2304 42400 2312 42464
rect 1992 41376 2312 42400
rect 1992 41312 2000 41376
rect 2064 41312 2080 41376
rect 2144 41312 2160 41376
rect 2224 41312 2240 41376
rect 2304 41312 2312 41376
rect 1992 40288 2312 41312
rect 1992 40224 2000 40288
rect 2064 40224 2080 40288
rect 2144 40224 2160 40288
rect 2224 40224 2240 40288
rect 2304 40224 2312 40288
rect 1992 39200 2312 40224
rect 1992 39136 2000 39200
rect 2064 39136 2080 39200
rect 2144 39136 2160 39200
rect 2224 39136 2240 39200
rect 2304 39136 2312 39200
rect 1992 38112 2312 39136
rect 1992 38048 2000 38112
rect 2064 38048 2080 38112
rect 2144 38048 2160 38112
rect 2224 38048 2240 38112
rect 2304 38048 2312 38112
rect 1992 37024 2312 38048
rect 1992 36960 2000 37024
rect 2064 36960 2080 37024
rect 2144 36960 2160 37024
rect 2224 36960 2240 37024
rect 2304 36960 2312 37024
rect 400 35492 748 35514
rect 400 35428 422 35492
rect 486 35428 502 35492
rect 566 35428 582 35492
rect 646 35428 662 35492
rect 726 35428 748 35492
rect 400 35412 748 35428
rect 400 35348 422 35412
rect 486 35348 502 35412
rect 566 35348 582 35412
rect 646 35348 662 35412
rect 726 35348 748 35412
rect 400 35332 748 35348
rect 400 35268 422 35332
rect 486 35268 502 35332
rect 566 35268 582 35332
rect 646 35268 662 35332
rect 726 35268 748 35332
rect 400 35252 748 35268
rect 400 35188 422 35252
rect 486 35188 502 35252
rect 566 35188 582 35252
rect 646 35188 662 35252
rect 726 35188 748 35252
rect 400 35166 748 35188
rect 1992 35492 2312 36960
rect 1992 35428 2000 35492
rect 2064 35428 2080 35492
rect 2144 35428 2160 35492
rect 2224 35428 2240 35492
rect 2304 35428 2312 35492
rect 1992 35412 2312 35428
rect 1992 35348 2000 35412
rect 2064 35348 2080 35412
rect 2144 35348 2160 35412
rect 2224 35348 2240 35412
rect 2304 35348 2312 35412
rect 1992 35332 2312 35348
rect 1992 35268 2000 35332
rect 2064 35268 2080 35332
rect 2144 35268 2160 35332
rect 2224 35268 2240 35332
rect 2304 35268 2312 35332
rect 1992 35252 2312 35268
rect 1992 35188 2000 35252
rect 2064 35188 2080 35252
rect 2144 35188 2160 35252
rect 2224 35188 2240 35252
rect 2304 35188 2312 35252
rect 1096 34796 1444 34818
rect 1096 34732 1118 34796
rect 1182 34732 1198 34796
rect 1262 34732 1278 34796
rect 1342 34732 1358 34796
rect 1422 34732 1444 34796
rect 1096 34716 1444 34732
rect 1096 34652 1118 34716
rect 1182 34652 1198 34716
rect 1262 34652 1278 34716
rect 1342 34652 1358 34716
rect 1422 34652 1444 34716
rect 1096 34636 1444 34652
rect 1096 34572 1118 34636
rect 1182 34572 1198 34636
rect 1262 34572 1278 34636
rect 1342 34572 1358 34636
rect 1422 34572 1444 34636
rect 1096 34556 1444 34572
rect 1096 34492 1118 34556
rect 1182 34492 1198 34556
rect 1262 34492 1278 34556
rect 1342 34492 1358 34556
rect 1422 34492 1444 34556
rect 1096 34470 1444 34492
rect 1992 34208 2312 35188
rect 2912 44096 3232 44656
rect 6134 44573 6194 45152
rect 6686 44573 6746 45152
rect 7238 44573 7298 45152
rect 7790 44573 7850 45152
rect 8342 44573 8402 45152
rect 8894 44573 8954 45152
rect 9446 44573 9506 45152
rect 9998 44573 10058 45152
rect 10550 44573 10610 45152
rect 11102 44573 11162 45152
rect 11654 44709 11714 45152
rect 11651 44708 11717 44709
rect 11651 44644 11652 44708
rect 11716 44644 11717 44708
rect 11651 44643 11717 44644
rect 12206 44573 12266 45152
rect 6131 44572 6197 44573
rect 6131 44508 6132 44572
rect 6196 44508 6197 44572
rect 6131 44507 6197 44508
rect 6683 44572 6749 44573
rect 6683 44508 6684 44572
rect 6748 44508 6749 44572
rect 6683 44507 6749 44508
rect 7235 44572 7301 44573
rect 7235 44508 7236 44572
rect 7300 44508 7301 44572
rect 7235 44507 7301 44508
rect 7787 44572 7853 44573
rect 7787 44508 7788 44572
rect 7852 44508 7853 44572
rect 7787 44507 7853 44508
rect 8339 44572 8405 44573
rect 8339 44508 8340 44572
rect 8404 44508 8405 44572
rect 8339 44507 8405 44508
rect 8891 44572 8957 44573
rect 8891 44508 8892 44572
rect 8956 44508 8957 44572
rect 8891 44507 8957 44508
rect 9443 44572 9509 44573
rect 9443 44508 9444 44572
rect 9508 44508 9509 44572
rect 9443 44507 9509 44508
rect 9995 44572 10061 44573
rect 9995 44508 9996 44572
rect 10060 44508 10061 44572
rect 9995 44507 10061 44508
rect 10547 44572 10613 44573
rect 10547 44508 10548 44572
rect 10612 44508 10613 44572
rect 10547 44507 10613 44508
rect 11099 44572 11165 44573
rect 11099 44508 11100 44572
rect 11164 44508 11165 44572
rect 11099 44507 11165 44508
rect 12203 44572 12269 44573
rect 12203 44508 12204 44572
rect 12268 44508 12269 44572
rect 12203 44507 12269 44508
rect 2912 44032 2920 44096
rect 2984 44032 3000 44096
rect 3064 44032 3080 44096
rect 3144 44032 3160 44096
rect 3224 44032 3232 44096
rect 2912 43008 3232 44032
rect 12758 43893 12818 45152
rect 13310 44845 13370 45152
rect 13862 44845 13922 45152
rect 13307 44844 13373 44845
rect 13307 44780 13308 44844
rect 13372 44780 13373 44844
rect 13307 44779 13373 44780
rect 13859 44844 13925 44845
rect 13859 44780 13860 44844
rect 13924 44780 13925 44844
rect 13859 44779 13925 44780
rect 14414 44573 14474 45152
rect 14966 44709 15026 45152
rect 14963 44708 15029 44709
rect 14963 44644 14964 44708
rect 15028 44644 15029 44708
rect 14963 44643 15029 44644
rect 15518 44573 15578 45152
rect 14411 44572 14477 44573
rect 14411 44508 14412 44572
rect 14476 44508 14477 44572
rect 14411 44507 14477 44508
rect 15515 44572 15581 44573
rect 15515 44508 15516 44572
rect 15580 44508 15581 44572
rect 15515 44507 15581 44508
rect 16070 43893 16130 45152
rect 12755 43892 12821 43893
rect 12755 43828 12756 43892
rect 12820 43828 12821 43892
rect 12755 43827 12821 43828
rect 16067 43892 16133 43893
rect 16067 43828 16068 43892
rect 16132 43828 16133 43892
rect 16067 43827 16133 43828
rect 2912 42944 2920 43008
rect 2984 42944 3000 43008
rect 3064 42944 3080 43008
rect 3144 42944 3160 43008
rect 3224 42944 3232 43008
rect 2912 41920 3232 42944
rect 16622 42941 16682 45152
rect 17174 43485 17234 45152
rect 17726 44573 17786 45152
rect 17723 44572 17789 44573
rect 17723 44508 17724 44572
rect 17788 44508 17789 44572
rect 17723 44507 17789 44508
rect 18278 44029 18338 45152
rect 18275 44028 18341 44029
rect 18275 43964 18276 44028
rect 18340 43964 18341 44028
rect 18275 43963 18341 43964
rect 17171 43484 17237 43485
rect 17171 43420 17172 43484
rect 17236 43420 17237 43484
rect 17171 43419 17237 43420
rect 16619 42940 16685 42941
rect 16619 42876 16620 42940
rect 16684 42876 16685 42940
rect 16619 42875 16685 42876
rect 18830 42397 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 18827 42396 18893 42397
rect 18827 42332 18828 42396
rect 18892 42332 18893 42396
rect 18827 42331 18893 42332
rect 2912 41856 2920 41920
rect 2984 41856 3000 41920
rect 3064 41856 3080 41920
rect 3144 41856 3160 41920
rect 3224 41856 3232 41920
rect 2912 40832 3232 41856
rect 2912 40768 2920 40832
rect 2984 40768 3000 40832
rect 3064 40768 3080 40832
rect 3144 40768 3160 40832
rect 3224 40768 3232 40832
rect 2912 39744 3232 40768
rect 3923 40628 3989 40629
rect 3923 40564 3924 40628
rect 3988 40564 3989 40628
rect 3923 40563 3989 40564
rect 2912 39680 2920 39744
rect 2984 39680 3000 39744
rect 3064 39680 3080 39744
rect 3144 39680 3160 39744
rect 3224 39680 3232 39744
rect 2912 38656 3232 39680
rect 2912 38592 2920 38656
rect 2984 38592 3000 38656
rect 3064 38592 3080 38656
rect 3144 38592 3160 38656
rect 3224 38592 3232 38656
rect 2912 37568 3232 38592
rect 2912 37504 2920 37568
rect 2984 37504 3000 37568
rect 3064 37504 3080 37568
rect 3144 37504 3160 37568
rect 3224 37504 3232 37568
rect 2912 34796 3232 37504
rect 3926 35910 3986 40563
rect 15515 39812 15581 39813
rect 15515 39748 15516 39812
rect 15580 39748 15581 39812
rect 15515 39747 15581 39748
rect 14411 37228 14477 37229
rect 14411 37164 14412 37228
rect 14476 37164 14477 37228
rect 14411 37163 14477 37164
rect 12019 37092 12085 37093
rect 12019 37028 12020 37092
rect 12084 37028 12085 37092
rect 12019 37027 12085 37028
rect 10915 36956 10981 36957
rect 10915 36892 10916 36956
rect 10980 36892 10981 36956
rect 10915 36891 10981 36892
rect 9627 36820 9693 36821
rect 9627 36756 9628 36820
rect 9692 36756 9693 36820
rect 9627 36755 9693 36756
rect 5027 36684 5093 36685
rect 5027 36620 5028 36684
rect 5092 36620 5093 36684
rect 5027 36619 5093 36620
rect 5030 35910 5090 36619
rect 6131 36548 6197 36549
rect 6131 36484 6132 36548
rect 6196 36484 6197 36548
rect 6131 36483 6197 36484
rect 3834 35850 3986 35910
rect 4984 35850 5090 35910
rect 3834 35476 3894 35850
rect 4984 35476 5044 35850
rect 6134 35476 6194 36483
rect 9630 35910 9690 36755
rect 10918 35910 10978 36891
rect 12022 35910 12082 37027
rect 13157 36004 13223 36005
rect 13157 35940 13158 36004
rect 13222 35940 13223 36004
rect 13157 35939 13223 35940
rect 9630 35850 9716 35910
rect 7327 35732 7393 35733
rect 7327 35668 7328 35732
rect 7392 35668 7393 35732
rect 7327 35667 7393 35668
rect 8485 35732 8551 35733
rect 8485 35668 8486 35732
rect 8550 35668 8551 35732
rect 8485 35667 8551 35668
rect 7330 35476 7390 35667
rect 8488 35476 8548 35667
rect 9656 35476 9716 35850
rect 10826 35850 10978 35910
rect 11992 35850 12082 35910
rect 10826 35476 10886 35850
rect 11992 35476 12052 35850
rect 13160 35476 13220 35939
rect 14414 35910 14474 37163
rect 15518 35910 15578 39747
rect 19011 39404 19077 39405
rect 19011 39340 19012 39404
rect 19076 39340 19077 39404
rect 19011 39339 19077 39340
rect 16619 36140 16685 36141
rect 16619 36076 16620 36140
rect 16684 36076 16685 36140
rect 16619 36075 16685 36076
rect 14322 35850 14474 35910
rect 15496 35850 15578 35910
rect 16622 35910 16682 36075
rect 16622 35850 16724 35910
rect 14322 35476 14382 35850
rect 15496 35476 15556 35850
rect 16664 35476 16724 35850
rect 17829 35868 17895 35869
rect 17829 35804 17830 35868
rect 17894 35804 17895 35868
rect 17829 35803 17895 35804
rect 17832 35476 17892 35803
rect 19014 35476 19074 39339
rect 21403 38316 21469 38317
rect 21403 38252 21404 38316
rect 21468 38252 21469 38316
rect 21403 38251 21469 38252
rect 20115 38044 20181 38045
rect 20115 37980 20116 38044
rect 20180 37980 20181 38044
rect 20115 37979 20181 37980
rect 20118 35910 20178 37979
rect 21406 35910 21466 38251
rect 21590 36277 21650 45152
rect 22142 43349 22202 45152
rect 22139 43348 22205 43349
rect 22139 43284 22140 43348
rect 22204 43284 22205 43348
rect 22139 43283 22205 43284
rect 22694 37229 22754 45152
rect 23246 43485 23306 45152
rect 23243 43484 23309 43485
rect 23243 43420 23244 43484
rect 23308 43420 23309 43484
rect 23243 43419 23309 43420
rect 23798 40629 23858 45152
rect 24350 41430 24410 45152
rect 24715 43348 24781 43349
rect 24715 43284 24716 43348
rect 24780 43284 24781 43348
rect 24715 43283 24781 43284
rect 24350 41370 24594 41430
rect 23795 40628 23861 40629
rect 23795 40564 23796 40628
rect 23860 40564 23861 40628
rect 23795 40563 23861 40564
rect 24347 40084 24413 40085
rect 24347 40020 24348 40084
rect 24412 40020 24413 40084
rect 24347 40019 24413 40020
rect 22691 37228 22757 37229
rect 22691 37164 22692 37228
rect 22756 37164 22757 37228
rect 22691 37163 22757 37164
rect 23611 37092 23677 37093
rect 23611 37028 23612 37092
rect 23676 37028 23677 37092
rect 23611 37027 23677 37028
rect 22507 36412 22573 36413
rect 22507 36348 22508 36412
rect 22572 36348 22573 36412
rect 22507 36347 22573 36348
rect 21587 36276 21653 36277
rect 21587 36212 21588 36276
rect 21652 36212 21653 36276
rect 21587 36211 21653 36212
rect 19471 35868 19537 35869
rect 19471 35804 19472 35868
rect 19536 35804 19537 35868
rect 20118 35850 20228 35910
rect 19471 35803 19537 35804
rect 19474 35476 19534 35803
rect 20027 35732 20093 35733
rect 20027 35668 20028 35732
rect 20092 35668 20093 35732
rect 20027 35667 20093 35668
rect 20030 35476 20090 35667
rect 20168 35476 20228 35850
rect 20967 35868 21033 35869
rect 20967 35804 20968 35868
rect 21032 35804 21033 35868
rect 20967 35803 21033 35804
rect 21336 35850 21466 35910
rect 20970 35476 21030 35803
rect 21195 35732 21261 35733
rect 21195 35668 21196 35732
rect 21260 35668 21261 35732
rect 21195 35667 21261 35668
rect 21198 35476 21258 35667
rect 21336 35476 21396 35850
rect 21967 35732 22033 35733
rect 21967 35668 21968 35732
rect 22032 35668 22033 35732
rect 21967 35667 22033 35668
rect 22139 35732 22205 35733
rect 22139 35668 22140 35732
rect 22204 35730 22205 35732
rect 22204 35668 22260 35730
rect 22139 35667 22260 35668
rect 21970 35476 22030 35667
rect 22200 35476 22260 35667
rect 22510 35476 22570 36347
rect 23614 36002 23674 37027
rect 23614 35942 23732 36002
rect 23197 35868 23263 35869
rect 23197 35804 23198 35868
rect 23262 35804 23263 35868
rect 23197 35803 23263 35804
rect 22967 35732 23033 35733
rect 22967 35668 22968 35732
rect 23032 35668 23033 35732
rect 22967 35667 23033 35668
rect 22970 35476 23030 35667
rect 23200 35476 23260 35803
rect 23531 35732 23597 35733
rect 23531 35668 23532 35732
rect 23596 35668 23597 35732
rect 23531 35667 23597 35668
rect 23534 35476 23594 35667
rect 23672 35476 23732 35942
rect 24350 35730 24410 40019
rect 24534 38589 24594 41370
rect 24531 38588 24597 38589
rect 24531 38524 24532 38588
rect 24596 38524 24597 38588
rect 24531 38523 24597 38524
rect 24718 37365 24778 43283
rect 24902 42941 24962 45152
rect 24899 42940 24965 42941
rect 24899 42876 24900 42940
rect 24964 42876 24965 42940
rect 24899 42875 24965 42876
rect 25454 40629 25514 45152
rect 26006 44981 26066 45152
rect 26003 44980 26069 44981
rect 26003 44916 26004 44980
rect 26068 44916 26069 44980
rect 26003 44915 26069 44916
rect 26558 44437 26618 45152
rect 27110 44709 27170 45152
rect 27662 44845 27722 45152
rect 27659 44844 27725 44845
rect 27659 44780 27660 44844
rect 27724 44780 27725 44844
rect 27659 44779 27725 44780
rect 28214 44709 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 27107 44708 27173 44709
rect 27107 44644 27108 44708
rect 27172 44644 27173 44708
rect 27107 44643 27173 44644
rect 28211 44708 28277 44709
rect 28211 44644 28212 44708
rect 28276 44644 28277 44708
rect 28211 44643 28277 44644
rect 49992 44640 50312 44656
rect 49992 44576 50000 44640
rect 50064 44576 50080 44640
rect 50144 44576 50160 44640
rect 50224 44576 50240 44640
rect 50304 44576 50312 44640
rect 26555 44436 26621 44437
rect 26555 44372 26556 44436
rect 26620 44372 26621 44436
rect 26555 44371 26621 44372
rect 49992 43552 50312 44576
rect 49992 43488 50000 43552
rect 50064 43488 50080 43552
rect 50144 43488 50160 43552
rect 50224 43488 50240 43552
rect 50304 43488 50312 43552
rect 32075 43484 32141 43485
rect 32075 43420 32076 43484
rect 32140 43420 32141 43484
rect 32075 43419 32141 43420
rect 27475 43076 27541 43077
rect 27475 43012 27476 43076
rect 27540 43012 27541 43076
rect 27475 43011 27541 43012
rect 27659 43076 27725 43077
rect 27659 43012 27660 43076
rect 27724 43012 27725 43076
rect 27659 43011 27725 43012
rect 26923 41036 26989 41037
rect 26923 40972 26924 41036
rect 26988 40972 26989 41036
rect 26923 40971 26989 40972
rect 25451 40628 25517 40629
rect 25451 40564 25452 40628
rect 25516 40564 25517 40628
rect 25451 40563 25517 40564
rect 26187 38724 26253 38725
rect 26187 38660 26188 38724
rect 26252 38660 26253 38724
rect 26187 38659 26253 38660
rect 26003 38452 26069 38453
rect 26003 38388 26004 38452
rect 26068 38388 26069 38452
rect 26003 38387 26069 38388
rect 24715 37364 24781 37365
rect 24715 37300 24716 37364
rect 24780 37300 24781 37364
rect 24715 37299 24781 37300
rect 24899 37228 24965 37229
rect 24899 37164 24900 37228
rect 24964 37164 24965 37228
rect 24899 37163 24965 37164
rect 24691 36004 24757 36005
rect 24691 35940 24692 36004
rect 24756 35940 24757 36004
rect 24902 36002 24962 37163
rect 24691 35939 24757 35940
rect 24840 35942 24962 36002
rect 24350 35670 24536 35730
rect 24476 35476 24536 35670
rect 24694 35476 24754 35939
rect 24840 35476 24900 35942
rect 25867 35868 25933 35869
rect 25867 35804 25868 35868
rect 25932 35804 25933 35868
rect 25867 35803 25933 35804
rect 25209 35732 25275 35733
rect 25209 35668 25210 35732
rect 25274 35668 25275 35732
rect 25209 35667 25275 35668
rect 25212 35476 25272 35667
rect 25870 35476 25930 35803
rect 26006 35476 26066 38387
rect 26190 35733 26250 38659
rect 26739 36548 26805 36549
rect 26739 36484 26740 36548
rect 26804 36484 26805 36548
rect 26739 36483 26805 36484
rect 26463 36004 26529 36005
rect 26463 35940 26464 36004
rect 26528 35940 26529 36004
rect 26742 36002 26802 36483
rect 26463 35939 26529 35940
rect 26694 35942 26802 36002
rect 26187 35732 26253 35733
rect 26187 35668 26188 35732
rect 26252 35668 26253 35732
rect 26187 35667 26253 35668
rect 26466 35476 26526 35939
rect 26694 35476 26754 35942
rect 26926 35730 26986 40971
rect 27478 40765 27538 43011
rect 27475 40764 27541 40765
rect 27475 40700 27476 40764
rect 27540 40700 27541 40764
rect 27475 40699 27541 40700
rect 27291 37500 27357 37501
rect 27291 37436 27292 37500
rect 27356 37436 27357 37500
rect 27291 37435 27357 37436
rect 27294 35910 27354 37435
rect 27662 36002 27722 43011
rect 30971 42124 31037 42125
rect 30971 42060 30972 42124
rect 31036 42060 31037 42124
rect 30971 42059 31037 42060
rect 27843 40356 27909 40357
rect 27843 40292 27844 40356
rect 27908 40292 27909 40356
rect 27843 40291 27909 40292
rect 27846 39269 27906 40291
rect 28579 39948 28645 39949
rect 28579 39884 28580 39948
rect 28644 39884 28645 39948
rect 28579 39883 28645 39884
rect 27843 39268 27909 39269
rect 27843 39204 27844 39268
rect 27908 39204 27909 39268
rect 27843 39203 27909 39204
rect 28395 38724 28461 38725
rect 28395 38660 28396 38724
rect 28460 38660 28461 38724
rect 28395 38659 28461 38660
rect 28027 37908 28093 37909
rect 28027 37844 28028 37908
rect 28092 37844 28093 37908
rect 28027 37843 28093 37844
rect 28030 37498 28090 37843
rect 27846 37438 28090 37498
rect 27846 37365 27906 37438
rect 27843 37364 27909 37365
rect 27843 37300 27844 37364
rect 27908 37300 27909 37364
rect 27843 37299 27909 37300
rect 28211 37228 28277 37229
rect 28211 37164 28212 37228
rect 28276 37164 28277 37228
rect 28211 37163 28277 37164
rect 27662 35942 27754 36002
rect 27176 35850 27354 35910
rect 26926 35670 27078 35730
rect 27018 35476 27078 35670
rect 27176 35476 27236 35850
rect 27694 35476 27754 35942
rect 28214 35476 28274 37163
rect 28398 36002 28458 38659
rect 28582 37501 28642 39883
rect 28947 38996 29013 38997
rect 28947 38932 28948 38996
rect 29012 38932 29013 38996
rect 28947 38931 29013 38932
rect 28579 37500 28645 37501
rect 28579 37436 28580 37500
rect 28644 37436 28645 37500
rect 28579 37435 28645 37436
rect 28344 35942 28458 36002
rect 28344 35476 28404 35942
rect 28950 35476 29010 38931
rect 29197 36004 29263 36005
rect 29197 35940 29198 36004
rect 29262 35940 29263 36004
rect 29197 35939 29263 35940
rect 30677 36004 30743 36005
rect 30677 35940 30678 36004
rect 30742 35940 30743 36004
rect 30974 36002 31034 42059
rect 31891 37500 31957 37501
rect 31891 37436 31892 37500
rect 31956 37436 31957 37500
rect 31891 37435 31957 37436
rect 31197 36004 31263 36005
rect 30974 35942 31101 36002
rect 30677 35939 30743 35940
rect 29200 35476 29260 35939
rect 29509 35868 29575 35869
rect 29509 35804 29510 35868
rect 29574 35804 29575 35868
rect 29509 35803 29575 35804
rect 30235 35868 30301 35869
rect 30235 35804 30236 35868
rect 30300 35804 30301 35868
rect 30235 35803 30301 35804
rect 29512 35476 29572 35803
rect 29967 35732 30033 35733
rect 29967 35668 29968 35732
rect 30032 35668 30033 35732
rect 30238 35730 30298 35803
rect 29967 35667 30033 35668
rect 30200 35670 30298 35730
rect 29970 35476 30030 35667
rect 30200 35476 30260 35670
rect 30680 35476 30740 35939
rect 31041 35476 31101 35942
rect 31197 35940 31198 36004
rect 31262 35940 31263 36004
rect 31197 35939 31263 35940
rect 31707 36004 31773 36005
rect 31707 35940 31708 36004
rect 31772 35940 31773 36004
rect 31707 35939 31773 35940
rect 31200 35476 31260 35939
rect 31710 35476 31770 35939
rect 31894 35910 31954 37435
rect 32078 36005 32138 43419
rect 35203 43212 35269 43213
rect 35203 43148 35204 43212
rect 35268 43148 35269 43212
rect 35203 43147 35269 43148
rect 35019 41308 35085 41309
rect 35019 41244 35020 41308
rect 35084 41244 35085 41308
rect 35019 41243 35085 41244
rect 32995 40900 33061 40901
rect 32995 40836 32996 40900
rect 33060 40836 33061 40900
rect 32995 40835 33061 40836
rect 32811 40628 32877 40629
rect 32811 40564 32812 40628
rect 32876 40564 32877 40628
rect 32811 40563 32877 40564
rect 32814 39269 32874 40563
rect 32998 39677 33058 40835
rect 32995 39676 33061 39677
rect 32995 39612 32996 39676
rect 33060 39612 33061 39676
rect 32995 39611 33061 39612
rect 32811 39268 32877 39269
rect 32811 39204 32812 39268
rect 32876 39204 32877 39268
rect 32811 39203 32877 39204
rect 32443 38724 32509 38725
rect 32443 38660 32444 38724
rect 32508 38660 32509 38724
rect 32443 38659 32509 38660
rect 33179 38724 33245 38725
rect 33179 38660 33180 38724
rect 33244 38660 33245 38724
rect 33179 38659 33245 38660
rect 32075 36004 32141 36005
rect 32075 35940 32076 36004
rect 32140 35940 32141 36004
rect 32075 35939 32141 35940
rect 31848 35850 31954 35910
rect 32446 35910 32506 38659
rect 32995 37500 33061 37501
rect 32995 37436 32996 37500
rect 33060 37436 33061 37500
rect 32995 37435 33061 37436
rect 32998 35910 33058 37435
rect 33182 36413 33242 38659
rect 34099 38588 34165 38589
rect 34099 38524 34100 38588
rect 34164 38524 34165 38588
rect 34099 38523 34165 38524
rect 33179 36412 33245 36413
rect 33179 36348 33180 36412
rect 33244 36348 33245 36412
rect 33179 36347 33245 36348
rect 34102 35910 34162 38523
rect 35022 35910 35082 41243
rect 32446 35850 32536 35910
rect 32998 35850 33076 35910
rect 31848 35476 31908 35850
rect 32476 35476 32536 35850
rect 32875 35732 32941 35733
rect 32875 35668 32876 35732
rect 32940 35668 32941 35732
rect 32875 35667 32941 35668
rect 32878 35476 32938 35667
rect 33016 35476 33076 35850
rect 33915 35868 33981 35869
rect 33915 35804 33916 35868
rect 33980 35804 33981 35868
rect 34102 35850 34254 35910
rect 33915 35803 33981 35804
rect 33455 35732 33521 35733
rect 33455 35668 33456 35732
rect 33520 35668 33521 35732
rect 33731 35732 33797 35733
rect 33731 35730 33732 35732
rect 33455 35667 33521 35668
rect 33694 35668 33732 35730
rect 33796 35668 33797 35732
rect 33918 35730 33978 35803
rect 33918 35670 34106 35730
rect 33694 35667 33797 35668
rect 33458 35476 33518 35667
rect 33694 35476 33754 35667
rect 34046 35476 34106 35670
rect 34194 35476 34254 35850
rect 34970 35850 35082 35910
rect 34970 35476 35030 35850
rect 35206 35476 35266 43147
rect 49992 42464 50312 43488
rect 49992 42400 50000 42464
rect 50064 42400 50080 42464
rect 50144 42400 50160 42464
rect 50224 42400 50240 42464
rect 50304 42400 50312 42464
rect 49992 41376 50312 42400
rect 49992 41312 50000 41376
rect 50064 41312 50080 41376
rect 50144 41312 50160 41376
rect 50224 41312 50240 41376
rect 50304 41312 50312 41376
rect 49992 40288 50312 41312
rect 49992 40224 50000 40288
rect 50064 40224 50080 40288
rect 50144 40224 50160 40288
rect 50224 40224 50240 40288
rect 50304 40224 50312 40288
rect 36123 39676 36189 39677
rect 36123 39612 36124 39676
rect 36188 39612 36189 39676
rect 36123 39611 36189 39612
rect 35387 38724 35453 38725
rect 35387 38660 35388 38724
rect 35452 38660 35453 38724
rect 35387 38659 35453 38660
rect 35390 35910 35450 38659
rect 35352 35850 35450 35910
rect 36126 35910 36186 39611
rect 49992 39200 50312 40224
rect 49992 39136 50000 39200
rect 50064 39136 50080 39200
rect 50144 39136 50160 39200
rect 50224 39136 50240 39200
rect 50304 39136 50312 39200
rect 46979 38724 47045 38725
rect 46979 38660 46980 38724
rect 47044 38660 47045 38724
rect 46979 38659 47045 38660
rect 45875 37364 45941 37365
rect 45875 37300 45876 37364
rect 45940 37300 45941 37364
rect 45875 37299 45941 37300
rect 38883 36956 38949 36957
rect 38883 36892 38884 36956
rect 38948 36892 38949 36956
rect 38883 36891 38949 36892
rect 37595 36820 37661 36821
rect 37595 36756 37596 36820
rect 37660 36756 37661 36820
rect 37595 36755 37661 36756
rect 37598 35910 37658 36755
rect 38886 35910 38946 36891
rect 39987 36684 40053 36685
rect 39987 36620 39988 36684
rect 40052 36620 40053 36684
rect 39987 36619 40053 36620
rect 36126 35850 36278 35910
rect 35352 35476 35412 35850
rect 36218 35476 36278 35850
rect 36517 35868 36583 35869
rect 36517 35804 36518 35868
rect 36582 35804 36583 35868
rect 37598 35850 37750 35910
rect 36517 35803 36583 35804
rect 36520 35476 36580 35803
rect 37690 35476 37750 35850
rect 38856 35850 38946 35910
rect 39990 35910 40050 36619
rect 39990 35850 40084 35910
rect 38856 35476 38916 35850
rect 40024 35476 40084 35850
rect 42357 35868 42423 35869
rect 42357 35804 42358 35868
rect 42422 35804 42423 35868
rect 42357 35803 42423 35804
rect 43525 35868 43591 35869
rect 43525 35804 43526 35868
rect 43590 35804 43591 35868
rect 43525 35803 43591 35804
rect 41183 35732 41249 35733
rect 41183 35668 41184 35732
rect 41248 35668 41249 35732
rect 41183 35667 41249 35668
rect 41186 35476 41246 35667
rect 42360 35476 42420 35803
rect 43528 35476 43588 35803
rect 44679 35732 44745 35733
rect 44679 35668 44680 35732
rect 44744 35668 44745 35732
rect 44679 35667 44745 35668
rect 44682 35476 44742 35667
rect 45878 35476 45938 37299
rect 46982 35730 47042 38659
rect 49992 38112 50312 39136
rect 49992 38048 50000 38112
rect 50064 38048 50080 38112
rect 50144 38048 50160 38112
rect 50224 38048 50240 38112
rect 50304 38048 50312 38112
rect 49992 37024 50312 38048
rect 49992 36960 50000 37024
rect 50064 36960 50080 37024
rect 50144 36960 50160 37024
rect 50224 36960 50240 37024
rect 50304 36960 50312 37024
rect 46982 35670 47092 35730
rect 47032 35476 47092 35670
rect 49992 35492 50312 36960
rect 2912 34732 2920 34796
rect 2984 34732 3000 34796
rect 3064 34732 3080 34796
rect 3144 34732 3160 34796
rect 3224 34732 3232 34796
rect 2912 34716 3232 34732
rect 2912 34652 2920 34716
rect 2984 34652 3000 34716
rect 3064 34652 3080 34716
rect 3144 34652 3160 34716
rect 3224 34652 3232 34716
rect 2912 34636 3232 34652
rect 2912 34572 2920 34636
rect 2984 34572 3000 34636
rect 3064 34572 3080 34636
rect 3144 34572 3160 34636
rect 3224 34572 3232 34636
rect 2912 34556 3232 34572
rect 2912 34492 2920 34556
rect 2984 34492 3000 34556
rect 3064 34492 3080 34556
rect 3144 34492 3160 34556
rect 3224 34492 3232 34556
rect 2912 34210 3232 34492
rect 49992 35428 50000 35492
rect 50064 35428 50080 35492
rect 50144 35428 50160 35492
rect 50224 35428 50240 35492
rect 50304 35428 50312 35492
rect 49992 35412 50312 35428
rect 49992 35348 50000 35412
rect 50064 35348 50080 35412
rect 50144 35348 50160 35412
rect 50224 35348 50240 35412
rect 50304 35348 50312 35412
rect 49992 35332 50312 35348
rect 49992 35268 50000 35332
rect 50064 35268 50080 35332
rect 50144 35268 50160 35332
rect 50224 35268 50240 35332
rect 50304 35268 50312 35332
rect 49992 35252 50312 35268
rect 49992 35188 50000 35252
rect 50064 35188 50080 35252
rect 50144 35188 50160 35252
rect 50224 35188 50240 35252
rect 50304 35188 50312 35252
rect 49992 34142 50312 35188
rect 50912 44096 51232 44656
rect 50912 44032 50920 44096
rect 50984 44032 51000 44096
rect 51064 44032 51080 44096
rect 51144 44032 51160 44096
rect 51224 44032 51232 44096
rect 50912 43008 51232 44032
rect 50912 42944 50920 43008
rect 50984 42944 51000 43008
rect 51064 42944 51080 43008
rect 51144 42944 51160 43008
rect 51224 42944 51232 43008
rect 50912 41920 51232 42944
rect 50912 41856 50920 41920
rect 50984 41856 51000 41920
rect 51064 41856 51080 41920
rect 51144 41856 51160 41920
rect 51224 41856 51232 41920
rect 50912 40832 51232 41856
rect 50912 40768 50920 40832
rect 50984 40768 51000 40832
rect 51064 40768 51080 40832
rect 51144 40768 51160 40832
rect 51224 40768 51232 40832
rect 50912 39744 51232 40768
rect 50912 39680 50920 39744
rect 50984 39680 51000 39744
rect 51064 39680 51080 39744
rect 51144 39680 51160 39744
rect 51224 39680 51232 39744
rect 50912 38656 51232 39680
rect 50912 38592 50920 38656
rect 50984 38592 51000 38656
rect 51064 38592 51080 38656
rect 51144 38592 51160 38656
rect 51224 38592 51232 38656
rect 50912 37568 51232 38592
rect 62803 38588 62869 38589
rect 62803 38524 62804 38588
rect 62868 38524 62869 38588
rect 62803 38523 62869 38524
rect 50912 37504 50920 37568
rect 50984 37504 51000 37568
rect 51064 37504 51080 37568
rect 51144 37504 51160 37568
rect 51224 37504 51232 37568
rect 50912 34796 51232 37504
rect 62619 36820 62685 36821
rect 62619 36756 62620 36820
rect 62684 36756 62685 36820
rect 62619 36755 62685 36756
rect 56245 35732 56311 35733
rect 56245 35668 56246 35732
rect 56310 35668 56311 35732
rect 56245 35667 56311 35668
rect 56248 35476 56308 35667
rect 62188 35492 62536 35514
rect 62188 35428 62210 35492
rect 62274 35428 62290 35492
rect 62354 35428 62370 35492
rect 62434 35428 62450 35492
rect 62514 35428 62536 35492
rect 62188 35412 62536 35428
rect 62188 35348 62210 35412
rect 62274 35348 62290 35412
rect 62354 35348 62370 35412
rect 62434 35348 62450 35412
rect 62514 35348 62536 35412
rect 62188 35332 62536 35348
rect 62188 35268 62210 35332
rect 62274 35268 62290 35332
rect 62354 35268 62370 35332
rect 62434 35268 62450 35332
rect 62514 35268 62536 35332
rect 62188 35252 62536 35268
rect 62188 35188 62210 35252
rect 62274 35188 62290 35252
rect 62354 35188 62370 35252
rect 62434 35188 62450 35252
rect 62514 35188 62536 35252
rect 62188 35166 62536 35188
rect 50912 34732 50920 34796
rect 50984 34732 51000 34796
rect 51064 34732 51080 34796
rect 51144 34732 51160 34796
rect 51224 34732 51232 34796
rect 50912 34716 51232 34732
rect 50912 34652 50920 34716
rect 50984 34652 51000 34716
rect 51064 34652 51080 34716
rect 51144 34652 51160 34716
rect 51224 34652 51232 34716
rect 50912 34636 51232 34652
rect 50912 34572 50920 34636
rect 50984 34572 51000 34636
rect 51064 34572 51080 34636
rect 51144 34572 51160 34636
rect 51224 34572 51232 34636
rect 50912 34556 51232 34572
rect 50912 34492 50920 34556
rect 50984 34492 51000 34556
rect 51064 34492 51080 34556
rect 51144 34492 51160 34556
rect 51224 34492 51232 34556
rect 50912 34142 51232 34492
rect 61492 34796 61840 34818
rect 61492 34732 61514 34796
rect 61578 34732 61594 34796
rect 61658 34732 61674 34796
rect 61738 34732 61754 34796
rect 61818 34732 61840 34796
rect 61492 34716 61840 34732
rect 61492 34652 61514 34716
rect 61578 34652 61594 34716
rect 61658 34652 61674 34716
rect 61738 34652 61754 34716
rect 61818 34652 61840 34716
rect 61492 34636 61840 34652
rect 61492 34572 61514 34636
rect 61578 34572 61594 34636
rect 61658 34572 61674 34636
rect 61738 34572 61754 34636
rect 61818 34572 61840 34636
rect 61492 34556 61840 34572
rect 61492 34492 61514 34556
rect 61578 34492 61594 34556
rect 61658 34492 61674 34556
rect 61738 34492 61754 34556
rect 61818 34492 61840 34556
rect 61492 34470 61840 34492
rect 62622 15741 62682 36755
rect 62806 35597 62866 38523
rect 62987 37772 63053 37773
rect 62987 37708 62988 37772
rect 63052 37708 63053 37772
rect 62987 37707 63053 37708
rect 62803 35596 62869 35597
rect 62803 35532 62804 35596
rect 62868 35532 62869 35596
rect 62803 35531 62869 35532
rect 62990 26250 63050 37707
rect 64332 37024 64652 37584
rect 64332 36960 64340 37024
rect 64404 36960 64420 37024
rect 64484 36960 64500 37024
rect 64564 36960 64580 37024
rect 64644 36960 64652 37024
rect 64091 36004 64157 36005
rect 64091 35940 64092 36004
rect 64156 35940 64157 36004
rect 64091 35939 64157 35940
rect 63539 35868 63605 35869
rect 63539 35804 63540 35868
rect 63604 35804 63605 35868
rect 63539 35803 63605 35804
rect 62806 26190 63050 26250
rect 62806 17237 62866 26190
rect 62803 17236 62869 17237
rect 62803 17172 62804 17236
rect 62868 17172 62869 17236
rect 62803 17171 62869 17172
rect 62619 15740 62685 15741
rect 62619 15676 62620 15740
rect 62684 15676 62685 15740
rect 62619 15675 62685 15676
rect 63542 7445 63602 35803
rect 63723 35052 63789 35053
rect 63723 34988 63724 35052
rect 63788 34988 63789 35052
rect 63723 34987 63789 34988
rect 63726 17917 63786 34987
rect 63907 33148 63973 33149
rect 63907 33084 63908 33148
rect 63972 33084 63973 33148
rect 63907 33083 63973 33084
rect 63723 17916 63789 17917
rect 63723 17852 63724 17916
rect 63788 17852 63789 17916
rect 63723 17851 63789 17852
rect 63539 7444 63605 7445
rect 63539 7380 63540 7444
rect 63604 7380 63605 7444
rect 63539 7379 63605 7380
rect 63910 6901 63970 33083
rect 64094 32469 64154 35939
rect 64332 35936 64652 36960
rect 64332 35872 64340 35936
rect 64404 35872 64420 35936
rect 64484 35872 64500 35936
rect 64564 35872 64580 35936
rect 64644 35872 64652 35936
rect 64332 34848 64652 35872
rect 64332 34784 64340 34848
rect 64404 34784 64420 34848
rect 64484 34784 64500 34848
rect 64564 34784 64580 34848
rect 64644 34784 64652 34848
rect 64332 33760 64652 34784
rect 64332 33696 64340 33760
rect 64404 33696 64420 33760
rect 64484 33696 64500 33760
rect 64564 33696 64580 33760
rect 64644 33696 64652 33760
rect 64332 32672 64652 33696
rect 64332 32608 64340 32672
rect 64404 32608 64420 32672
rect 64484 32608 64500 32672
rect 64564 32608 64580 32672
rect 64644 32608 64652 32672
rect 64091 32468 64157 32469
rect 64091 32404 64092 32468
rect 64156 32404 64157 32468
rect 64091 32403 64157 32404
rect 64332 31584 64652 32608
rect 64332 31520 64340 31584
rect 64404 31520 64420 31584
rect 64484 31520 64500 31584
rect 64564 31520 64580 31584
rect 64644 31520 64652 31584
rect 64332 30496 64652 31520
rect 64332 30432 64340 30496
rect 64404 30432 64420 30496
rect 64484 30432 64500 30496
rect 64564 30432 64580 30496
rect 64644 30432 64652 30496
rect 64332 29408 64652 30432
rect 64332 29344 64340 29408
rect 64404 29344 64420 29408
rect 64484 29344 64500 29408
rect 64564 29344 64580 29408
rect 64644 29344 64652 29408
rect 64332 28320 64652 29344
rect 64332 28256 64340 28320
rect 64404 28256 64420 28320
rect 64484 28256 64500 28320
rect 64564 28256 64580 28320
rect 64644 28256 64652 28320
rect 64332 27232 64652 28256
rect 64332 27168 64340 27232
rect 64404 27168 64420 27232
rect 64484 27168 64500 27232
rect 64564 27168 64580 27232
rect 64644 27168 64652 27232
rect 64332 26144 64652 27168
rect 64332 26080 64340 26144
rect 64404 26080 64420 26144
rect 64484 26080 64500 26144
rect 64564 26080 64580 26144
rect 64644 26080 64652 26144
rect 64332 25056 64652 26080
rect 64332 24992 64340 25056
rect 64404 24992 64420 25056
rect 64484 24992 64500 25056
rect 64564 24992 64580 25056
rect 64644 24992 64652 25056
rect 64332 23968 64652 24992
rect 64332 23904 64340 23968
rect 64404 23904 64420 23968
rect 64484 23904 64500 23968
rect 64564 23904 64580 23968
rect 64644 23904 64652 23968
rect 64332 22880 64652 23904
rect 64332 22816 64340 22880
rect 64404 22816 64420 22880
rect 64484 22816 64500 22880
rect 64564 22816 64580 22880
rect 64644 22816 64652 22880
rect 64332 21792 64652 22816
rect 64332 21728 64340 21792
rect 64404 21728 64420 21792
rect 64484 21728 64500 21792
rect 64564 21728 64580 21792
rect 64644 21728 64652 21792
rect 64332 20704 64652 21728
rect 64332 20640 64340 20704
rect 64404 20640 64420 20704
rect 64484 20640 64500 20704
rect 64564 20640 64580 20704
rect 64644 20640 64652 20704
rect 64332 19616 64652 20640
rect 64332 19552 64340 19616
rect 64404 19552 64420 19616
rect 64484 19552 64500 19616
rect 64564 19552 64580 19616
rect 64644 19552 64652 19616
rect 64332 18528 64652 19552
rect 64332 18464 64340 18528
rect 64404 18464 64420 18528
rect 64484 18464 64500 18528
rect 64564 18464 64580 18528
rect 64644 18464 64652 18528
rect 64332 17440 64652 18464
rect 64332 17376 64340 17440
rect 64404 17376 64420 17440
rect 64484 17376 64500 17440
rect 64564 17376 64580 17440
rect 64644 17376 64652 17440
rect 64332 16352 64652 17376
rect 64332 16288 64340 16352
rect 64404 16288 64420 16352
rect 64484 16288 64500 16352
rect 64564 16288 64580 16352
rect 64644 16288 64652 16352
rect 64332 15264 64652 16288
rect 64332 15200 64340 15264
rect 64404 15200 64420 15264
rect 64484 15200 64500 15264
rect 64564 15200 64580 15264
rect 64644 15200 64652 15264
rect 64332 14176 64652 15200
rect 64332 14112 64340 14176
rect 64404 14112 64420 14176
rect 64484 14112 64500 14176
rect 64564 14112 64580 14176
rect 64644 14112 64652 14176
rect 64332 13088 64652 14112
rect 64332 13024 64340 13088
rect 64404 13024 64420 13088
rect 64484 13024 64500 13088
rect 64564 13024 64580 13088
rect 64644 13024 64652 13088
rect 64332 12000 64652 13024
rect 64332 11936 64340 12000
rect 64404 11936 64420 12000
rect 64484 11936 64500 12000
rect 64564 11936 64580 12000
rect 64644 11936 64652 12000
rect 64332 10912 64652 11936
rect 64332 10848 64340 10912
rect 64404 10848 64420 10912
rect 64484 10848 64500 10912
rect 64564 10848 64580 10912
rect 64644 10848 64652 10912
rect 64332 9824 64652 10848
rect 64332 9760 64340 9824
rect 64404 9760 64420 9824
rect 64484 9760 64500 9824
rect 64564 9760 64580 9824
rect 64644 9760 64652 9824
rect 64332 8736 64652 9760
rect 64332 8672 64340 8736
rect 64404 8672 64420 8736
rect 64484 8672 64500 8736
rect 64564 8672 64580 8736
rect 64644 8672 64652 8736
rect 64332 7648 64652 8672
rect 64332 7584 64340 7648
rect 64404 7584 64420 7648
rect 64484 7584 64500 7648
rect 64564 7584 64580 7648
rect 64644 7584 64652 7648
rect 63907 6900 63973 6901
rect 63907 6836 63908 6900
rect 63972 6836 63973 6900
rect 63907 6835 63973 6836
rect 64332 6560 64652 7584
rect 64332 6496 64340 6560
rect 64404 6496 64420 6560
rect 64484 6496 64500 6560
rect 64564 6496 64580 6560
rect 64644 6496 64652 6560
rect 64332 5472 64652 6496
rect 64332 5408 64340 5472
rect 64404 5408 64420 5472
rect 64484 5408 64500 5472
rect 64564 5408 64580 5472
rect 64644 5408 64652 5472
rect 64332 4384 64652 5408
rect 64332 4320 64340 4384
rect 64404 4320 64420 4384
rect 64484 4320 64500 4384
rect 64564 4320 64580 4384
rect 64644 4320 64652 4384
rect 64332 3296 64652 4320
rect 64332 3232 64340 3296
rect 64404 3232 64420 3296
rect 64484 3232 64500 3296
rect 64564 3232 64580 3296
rect 64644 3232 64652 3296
rect 1096 3022 1444 3044
rect 1096 2958 1118 3022
rect 1182 2958 1198 3022
rect 1262 2958 1278 3022
rect 1342 2958 1358 3022
rect 1422 2958 1444 3022
rect 1096 2942 1444 2958
rect 1096 2878 1118 2942
rect 1182 2878 1198 2942
rect 1262 2878 1278 2942
rect 1342 2878 1358 2942
rect 1422 2878 1444 2942
rect 1096 2862 1444 2878
rect 1096 2798 1118 2862
rect 1182 2798 1198 2862
rect 1262 2798 1278 2862
rect 1342 2798 1358 2862
rect 1422 2798 1444 2862
rect 1096 2782 1444 2798
rect 1096 2718 1118 2782
rect 1182 2718 1198 2782
rect 1262 2718 1278 2782
rect 1342 2718 1358 2782
rect 1422 2718 1444 2782
rect 1096 2696 1444 2718
rect 61492 3022 61840 3044
rect 61492 2958 61514 3022
rect 61578 2958 61594 3022
rect 61658 2958 61674 3022
rect 61738 2958 61754 3022
rect 61818 2958 61840 3022
rect 61492 2942 61840 2958
rect 61492 2878 61514 2942
rect 61578 2878 61594 2942
rect 61658 2878 61674 2942
rect 61738 2878 61754 2942
rect 61818 2878 61840 2942
rect 61492 2862 61840 2878
rect 61492 2798 61514 2862
rect 61578 2798 61594 2862
rect 61658 2798 61674 2862
rect 61738 2798 61754 2862
rect 61818 2798 61840 2862
rect 61492 2782 61840 2798
rect 61492 2718 61514 2782
rect 61578 2718 61594 2782
rect 61658 2718 61674 2782
rect 61738 2718 61754 2782
rect 61818 2718 61840 2782
rect 61492 2696 61840 2718
rect 400 2326 748 2348
rect 400 2262 422 2326
rect 486 2262 502 2326
rect 566 2262 582 2326
rect 646 2262 662 2326
rect 726 2262 748 2326
rect 400 2246 748 2262
rect 400 2182 422 2246
rect 486 2182 502 2246
rect 566 2182 582 2246
rect 646 2182 662 2246
rect 726 2182 748 2246
rect 400 2166 748 2182
rect 400 2102 422 2166
rect 486 2102 502 2166
rect 566 2102 582 2166
rect 646 2102 662 2166
rect 726 2102 748 2166
rect 400 2086 748 2102
rect 400 2022 422 2086
rect 486 2022 502 2086
rect 566 2022 582 2086
rect 646 2022 662 2086
rect 726 2022 748 2086
rect 62188 2326 62536 2348
rect 62188 2262 62210 2326
rect 62274 2262 62290 2326
rect 62354 2262 62370 2326
rect 62434 2262 62450 2326
rect 62514 2262 62536 2326
rect 62188 2246 62536 2262
rect 62188 2182 62210 2246
rect 62274 2182 62290 2246
rect 62354 2182 62370 2246
rect 62434 2182 62450 2246
rect 62514 2182 62536 2246
rect 62188 2166 62536 2182
rect 62188 2102 62210 2166
rect 62274 2102 62290 2166
rect 62354 2102 62370 2166
rect 62434 2102 62450 2166
rect 62514 2102 62536 2166
rect 62188 2086 62536 2102
rect 400 2000 748 2022
rect 48943 1869 49003 2038
rect 48940 1868 49006 1869
rect 48940 1804 48941 1868
rect 49005 1804 49006 1868
rect 48940 1803 49006 1804
rect 49081 1597 49141 2038
rect 49219 1597 49279 2038
rect 49374 1869 49434 2038
rect 49371 1868 49437 1869
rect 49371 1804 49372 1868
rect 49436 1804 49437 1868
rect 49371 1803 49437 1804
rect 49676 1733 49736 2038
rect 49673 1732 49739 1733
rect 49673 1668 49674 1732
rect 49738 1668 49739 1732
rect 49834 1730 49894 2038
rect 62188 2022 62210 2086
rect 62274 2022 62290 2086
rect 62354 2022 62370 2086
rect 62434 2022 62450 2086
rect 62514 2022 62536 2086
rect 62188 2000 62536 2022
rect 64332 2208 64652 3232
rect 64332 2144 64340 2208
rect 64404 2144 64420 2208
rect 64484 2144 64500 2208
rect 64564 2144 64580 2208
rect 64644 2144 64652 2208
rect 49834 1670 49986 1730
rect 49673 1667 49739 1668
rect 49078 1596 49144 1597
rect 49078 1532 49079 1596
rect 49143 1532 49144 1596
rect 49078 1531 49144 1532
rect 49216 1596 49282 1597
rect 49216 1532 49217 1596
rect 49281 1532 49282 1596
rect 49216 1531 49282 1532
rect 49926 1325 49986 1670
rect 49923 1324 49989 1325
rect 49923 1260 49924 1324
rect 49988 1260 49989 1324
rect 49923 1259 49989 1260
rect 64332 1120 64652 2144
rect 64332 1056 64340 1120
rect 64404 1056 64420 1120
rect 64484 1056 64500 1120
rect 64564 1056 64580 1120
rect 64644 1056 64652 1120
rect 64332 496 64652 1056
rect 65252 37568 65572 37584
rect 65252 37504 65260 37568
rect 65324 37504 65340 37568
rect 65404 37504 65420 37568
rect 65484 37504 65500 37568
rect 65564 37504 65572 37568
rect 65252 36480 65572 37504
rect 65252 36416 65260 36480
rect 65324 36416 65340 36480
rect 65404 36416 65420 36480
rect 65484 36416 65500 36480
rect 65564 36416 65572 36480
rect 65252 35392 65572 36416
rect 65252 35328 65260 35392
rect 65324 35328 65340 35392
rect 65404 35328 65420 35392
rect 65484 35328 65500 35392
rect 65564 35328 65572 35392
rect 65252 34304 65572 35328
rect 65252 34240 65260 34304
rect 65324 34240 65340 34304
rect 65404 34240 65420 34304
rect 65484 34240 65500 34304
rect 65564 34240 65572 34304
rect 65252 33216 65572 34240
rect 65252 33152 65260 33216
rect 65324 33152 65340 33216
rect 65404 33152 65420 33216
rect 65484 33152 65500 33216
rect 65564 33152 65572 33216
rect 65252 32128 65572 33152
rect 65252 32064 65260 32128
rect 65324 32064 65340 32128
rect 65404 32064 65420 32128
rect 65484 32064 65500 32128
rect 65564 32064 65572 32128
rect 65252 31040 65572 32064
rect 65252 30976 65260 31040
rect 65324 30976 65340 31040
rect 65404 30976 65420 31040
rect 65484 30976 65500 31040
rect 65564 30976 65572 31040
rect 65252 29952 65572 30976
rect 65252 29888 65260 29952
rect 65324 29888 65340 29952
rect 65404 29888 65420 29952
rect 65484 29888 65500 29952
rect 65564 29888 65572 29952
rect 65252 28864 65572 29888
rect 65252 28800 65260 28864
rect 65324 28800 65340 28864
rect 65404 28800 65420 28864
rect 65484 28800 65500 28864
rect 65564 28800 65572 28864
rect 65252 27776 65572 28800
rect 65252 27712 65260 27776
rect 65324 27712 65340 27776
rect 65404 27712 65420 27776
rect 65484 27712 65500 27776
rect 65564 27712 65572 27776
rect 65252 26688 65572 27712
rect 65252 26624 65260 26688
rect 65324 26624 65340 26688
rect 65404 26624 65420 26688
rect 65484 26624 65500 26688
rect 65564 26624 65572 26688
rect 65252 25600 65572 26624
rect 65252 25536 65260 25600
rect 65324 25536 65340 25600
rect 65404 25536 65420 25600
rect 65484 25536 65500 25600
rect 65564 25536 65572 25600
rect 65252 24512 65572 25536
rect 65252 24448 65260 24512
rect 65324 24448 65340 24512
rect 65404 24448 65420 24512
rect 65484 24448 65500 24512
rect 65564 24448 65572 24512
rect 65252 23424 65572 24448
rect 65252 23360 65260 23424
rect 65324 23360 65340 23424
rect 65404 23360 65420 23424
rect 65484 23360 65500 23424
rect 65564 23360 65572 23424
rect 65252 22336 65572 23360
rect 65252 22272 65260 22336
rect 65324 22272 65340 22336
rect 65404 22272 65420 22336
rect 65484 22272 65500 22336
rect 65564 22272 65572 22336
rect 65252 21248 65572 22272
rect 65252 21184 65260 21248
rect 65324 21184 65340 21248
rect 65404 21184 65420 21248
rect 65484 21184 65500 21248
rect 65564 21184 65572 21248
rect 65252 20160 65572 21184
rect 65252 20096 65260 20160
rect 65324 20096 65340 20160
rect 65404 20096 65420 20160
rect 65484 20096 65500 20160
rect 65564 20096 65572 20160
rect 65252 19072 65572 20096
rect 65252 19008 65260 19072
rect 65324 19008 65340 19072
rect 65404 19008 65420 19072
rect 65484 19008 65500 19072
rect 65564 19008 65572 19072
rect 65252 17984 65572 19008
rect 65252 17920 65260 17984
rect 65324 17920 65340 17984
rect 65404 17920 65420 17984
rect 65484 17920 65500 17984
rect 65564 17920 65572 17984
rect 65252 16896 65572 17920
rect 65252 16832 65260 16896
rect 65324 16832 65340 16896
rect 65404 16832 65420 16896
rect 65484 16832 65500 16896
rect 65564 16832 65572 16896
rect 65252 15808 65572 16832
rect 65252 15744 65260 15808
rect 65324 15744 65340 15808
rect 65404 15744 65420 15808
rect 65484 15744 65500 15808
rect 65564 15744 65572 15808
rect 65252 14720 65572 15744
rect 65252 14656 65260 14720
rect 65324 14656 65340 14720
rect 65404 14656 65420 14720
rect 65484 14656 65500 14720
rect 65564 14656 65572 14720
rect 65252 13632 65572 14656
rect 65252 13568 65260 13632
rect 65324 13568 65340 13632
rect 65404 13568 65420 13632
rect 65484 13568 65500 13632
rect 65564 13568 65572 13632
rect 65252 12544 65572 13568
rect 65252 12480 65260 12544
rect 65324 12480 65340 12544
rect 65404 12480 65420 12544
rect 65484 12480 65500 12544
rect 65564 12480 65572 12544
rect 65252 11456 65572 12480
rect 65252 11392 65260 11456
rect 65324 11392 65340 11456
rect 65404 11392 65420 11456
rect 65484 11392 65500 11456
rect 65564 11392 65572 11456
rect 65252 10368 65572 11392
rect 65252 10304 65260 10368
rect 65324 10304 65340 10368
rect 65404 10304 65420 10368
rect 65484 10304 65500 10368
rect 65564 10304 65572 10368
rect 65252 9280 65572 10304
rect 65252 9216 65260 9280
rect 65324 9216 65340 9280
rect 65404 9216 65420 9280
rect 65484 9216 65500 9280
rect 65564 9216 65572 9280
rect 65252 8192 65572 9216
rect 65252 8128 65260 8192
rect 65324 8128 65340 8192
rect 65404 8128 65420 8192
rect 65484 8128 65500 8192
rect 65564 8128 65572 8192
rect 65252 7104 65572 8128
rect 65252 7040 65260 7104
rect 65324 7040 65340 7104
rect 65404 7040 65420 7104
rect 65484 7040 65500 7104
rect 65564 7040 65572 7104
rect 65252 6016 65572 7040
rect 65252 5952 65260 6016
rect 65324 5952 65340 6016
rect 65404 5952 65420 6016
rect 65484 5952 65500 6016
rect 65564 5952 65572 6016
rect 65252 4928 65572 5952
rect 65252 4864 65260 4928
rect 65324 4864 65340 4928
rect 65404 4864 65420 4928
rect 65484 4864 65500 4928
rect 65564 4864 65572 4928
rect 65252 3840 65572 4864
rect 65252 3776 65260 3840
rect 65324 3776 65340 3840
rect 65404 3776 65420 3840
rect 65484 3776 65500 3840
rect 65564 3776 65572 3840
rect 65252 2752 65572 3776
rect 65252 2688 65260 2752
rect 65324 2688 65340 2752
rect 65404 2688 65420 2752
rect 65484 2688 65500 2752
rect 65564 2688 65572 2752
rect 65252 1664 65572 2688
rect 65252 1600 65260 1664
rect 65324 1600 65340 1664
rect 65404 1600 65420 1664
rect 65484 1600 65500 1664
rect 65564 1600 65572 1664
rect 65252 576 65572 1600
rect 65252 512 65260 576
rect 65324 512 65340 576
rect 65404 512 65420 576
rect 65484 512 65500 576
rect 65564 512 65572 576
rect 65252 496 65572 512
use sky130_fd_sc_hd__mux2_1  _250_
timestamp 1
transform -1 0 27416 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _251_
timestamp 1
transform 1 0 26680 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _252_
timestamp 1
transform -1 0 57592 0 1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _253_
timestamp 1
transform 1 0 12604 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _254_
timestamp 1
transform 1 0 10948 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _255_
timestamp 1
transform -1 0 8280 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _256_
timestamp 1
transform 1 0 10212 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _257_
timestamp 1
transform -1 0 22080 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _258_
timestamp 1
transform 1 0 22080 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _259_
timestamp 1
transform 1 0 9568 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _260_
timestamp 1
transform 1 0 9200 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _261_
timestamp 1
transform 1 0 8648 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _262_
timestamp 1
transform 1 0 9200 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _263_
timestamp 1
transform 1 0 10948 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _264_
timestamp 1
transform 1 0 7452 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _265_
timestamp 1
transform 1 0 9016 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _266_
timestamp 1
transform 1 0 12236 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _267_
timestamp 1
transform -1 0 10856 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _268_
timestamp 1
transform 1 0 11132 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _269_
timestamp 1
transform -1 0 60720 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _270_
timestamp 1
transform 1 0 59892 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _271_
timestamp 1
transform 1 0 58880 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _272_
timestamp 1
transform -1 0 57868 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _273_
timestamp 1
transform 1 0 58052 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _274_
timestamp 1
transform -1 0 57224 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _275_
timestamp 1
transform -1 0 56120 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _276_
timestamp 1
transform 1 0 55476 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _277_
timestamp 1
transform -1 0 56948 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _278_
timestamp 1
transform 1 0 54004 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _279_
timestamp 1
transform -1 0 53728 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _280_
timestamp 1
transform -1 0 54188 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _281_
timestamp 1
transform -1 0 55568 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _282_
timestamp 1
transform 1 0 54832 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _283_
timestamp 1
transform 1 0 55568 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _284_
timestamp 1
transform 1 0 52348 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _285_
timestamp 1
transform 1 0 52164 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _286_
timestamp 1
transform 1 0 53268 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _287_
timestamp 1
transform -1 0 20608 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _288_
timestamp 1
transform 1 0 22080 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _289_
timestamp 1
transform 1 0 52072 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _290_
timestamp 1
transform -1 0 50232 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _291_
timestamp 1
transform 1 0 49588 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _292_
timestamp 1
transform 1 0 50416 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _293_
timestamp 1
transform 1 0 48668 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _294_
timestamp 1
transform 1 0 48576 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _295_
timestamp 1
transform -1 0 50416 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _296_
timestamp 1
transform -1 0 48116 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _297_
timestamp 1
transform 1 0 48116 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _298_
timestamp 1
transform 1 0 47380 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _299_
timestamp 1
transform -1 0 47840 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _300_
timestamp 1
transform 1 0 47840 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _301_
timestamp 1
transform 1 0 47012 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _302_
timestamp 1
transform 1 0 45724 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _303_
timestamp 1
transform 1 0 45540 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _304_
timestamp 1
transform 1 0 45724 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _305_
timestamp 1
transform -1 0 46092 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _306_
timestamp 1
transform 1 0 46092 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _307_
timestamp 1
transform 1 0 45356 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _308_
timestamp 1
transform -1 0 45264 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _309_
timestamp 1
transform 1 0 44436 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _310_
timestamp 1
transform -1 0 46092 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _311_
timestamp 1
transform -1 0 42872 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _312_
timestamp 1
transform 1 0 42044 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _313_
timestamp 1
transform -1 0 43700 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _314_
timestamp 1
transform 1 0 41584 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _315_
timestamp 1
transform 1 0 40388 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _316_
timestamp 1
transform 1 0 42872 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _317_
timestamp 1
transform -1 0 17572 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _318_
timestamp 1
transform 1 0 18676 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _319_
timestamp 1
transform 1 0 39928 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _320_
timestamp 1
transform 1 0 39284 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _321_
timestamp 1
transform 1 0 38088 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _322_
timestamp 1
transform 1 0 39284 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _323_
timestamp 1
transform 1 0 35788 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _324_
timestamp 1
transform 1 0 34960 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _325_
timestamp 1
transform 1 0 36708 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _326_
timestamp 1
transform 1 0 33212 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _327_
timestamp 1
transform 1 0 32384 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _328_
timestamp 1
transform -1 0 34960 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _329_
timestamp 1
transform 1 0 31556 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _330_
timestamp 1
transform 1 0 30636 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _331_
timestamp 1
transform -1 0 31464 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _332_
timestamp 1
transform 1 0 30360 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _333_
timestamp 1
transform 1 0 29532 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _334_
timestamp 1
transform 1 0 30360 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _335_
timestamp 1
transform 1 0 28428 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _336_
timestamp 1
transform 1 0 28244 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _337_
timestamp 1
transform 1 0 29440 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _338_
timestamp 1
transform 1 0 27876 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _339_
timestamp 1
transform 1 0 27048 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _340_
timestamp 1
transform 1 0 27876 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _341_
timestamp 1
transform 1 0 26404 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _342_
timestamp 1
transform 1 0 25668 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _343_
timestamp 1
transform 1 0 25484 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _344_
timestamp 1
transform 1 0 25116 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _345_
timestamp 1
transform 1 0 23828 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _346_
timestamp 1
transform 1 0 25300 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _347_
timestamp 1
transform 1 0 17756 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _348_
timestamp 1
transform 1 0 15180 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _349_
timestamp 1
transform -1 0 24472 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _350_
timestamp 1
transform 1 0 21344 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _351_
timestamp 1
transform 1 0 19780 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1
transform 1 0 21252 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1
transform 1 0 18676 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _354_
timestamp 1
transform 1 0 17572 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _355_
timestamp 1
transform 1 0 18676 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _356_
timestamp 1
transform 1 0 16100 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _357_
timestamp 1
transform 1 0 14076 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _358_
timestamp 1
transform 1 0 15180 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _359_
timestamp 1
transform -1 0 14536 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _360_
timestamp 1
transform 1 0 13800 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _361_
timestamp 1
transform -1 0 13432 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _362_
timestamp 1
transform 1 0 12512 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _363_
timestamp 1
transform 1 0 11040 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _364_
timestamp 1
transform 1 0 11316 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _365_
timestamp 1
transform 1 0 15180 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _366_
timestamp 1
transform 1 0 14444 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _367_
timestamp 1
transform 1 0 13616 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _368_
timestamp 1
transform 1 0 43516 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _369_
timestamp 1
transform 1 0 41860 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _370_
timestamp 1
transform 1 0 44436 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _371_
timestamp 1
transform 1 0 40756 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _372_
timestamp 1
transform 1 0 43700 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _373_
timestamp 1
transform 1 0 41860 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _374_
timestamp 1
transform 1 0 43700 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _375_
timestamp 1
transform -1 0 41768 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _376_
timestamp 1
transform 1 0 44436 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _377_
timestamp 1
transform 1 0 43700 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _378_
timestamp 1
transform 1 0 43240 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _379_
timestamp 1
transform 1 0 42688 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1
transform 1 0 17296 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _381_
timestamp 1
transform 1 0 16468 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _382_
timestamp 1
transform -1 0 47840 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _383_
timestamp 1
transform -1 0 47840 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _384_
timestamp 1
transform 1 0 52164 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _385_
timestamp 1
transform 1 0 50876 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _386_
timestamp 1
transform 1 0 49956 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _387_
timestamp 1
transform 1 0 49864 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _388_
timestamp 1
transform 1 0 64676 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _389_
timestamp 1
transform 1 0 64216 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _390_
timestamp 1
transform -1 0 64676 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _391_
timestamp 1
transform 1 0 63848 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _392_
timestamp 1
transform 1 0 65320 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _393_
timestamp 1
transform 1 0 64584 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _394_
timestamp 1
transform -1 0 65320 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _395_
timestamp 1
transform 1 0 64584 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _396_
timestamp 1
transform -1 0 65412 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _397_
timestamp 1
transform 1 0 64860 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _398_
timestamp 1
transform 1 0 64676 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _399_
timestamp 1
transform 1 0 64492 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _400_
timestamp 1
transform 1 0 64584 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _401_
timestamp 1
transform 1 0 64584 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _402_
timestamp 1
transform -1 0 65320 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _403_
timestamp 1
transform 1 0 64584 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _404_
timestamp 1
transform 1 0 64584 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _405_
timestamp 1
transform 1 0 64584 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _406_
timestamp 1
transform -1 0 65412 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _407_
timestamp 1
transform 1 0 64584 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _408_
timestamp 1
transform 1 0 64584 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _409_
timestamp 1
transform 1 0 64584 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _410_
timestamp 1
transform -1 0 65320 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _411_
timestamp 1
transform 1 0 64584 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _412_
timestamp 1
transform -1 0 65412 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _413_
timestamp 1
transform 1 0 65320 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _414_
timestamp 1
transform -1 0 65228 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _415_
timestamp 1
transform 1 0 64492 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _416_
timestamp 1
transform 1 0 65044 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _417_
timestamp 1
transform 1 0 64676 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _418_
timestamp 1
transform -1 0 65136 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _419_
timestamp 1
transform 1 0 64492 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _420_
timestamp 1
transform -1 0 19872 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _421_
timestamp 1
transform 1 0 19228 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _422_
timestamp 1
transform -1 0 39192 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _423_
timestamp 1
transform 1 0 40112 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _424_
timestamp 1
transform -1 0 36616 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _425_
timestamp 1
transform 1 0 38548 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _426_
timestamp 1
transform 1 0 37628 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _427_
timestamp 1
transform 1 0 37260 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _428_
timestamp 1
transform -1 0 37536 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _429_
timestamp 1
transform 1 0 37812 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _430_
timestamp 1
transform 1 0 36708 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _431_
timestamp 1
transform 1 0 35788 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _432_
timestamp 1
transform -1 0 36616 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _433_
timestamp 1
transform -1 0 37536 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _434_
timestamp 1
transform -1 0 36616 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _435_
timestamp 1
transform 1 0 38180 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _436_
timestamp 1
transform 1 0 34960 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _437_
timestamp 1
transform 1 0 33212 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _438_
timestamp 1
transform -1 0 34868 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _439_
timestamp 1
transform 1 0 34132 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _440_
timestamp 1
transform 1 0 33212 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _441_
timestamp 1
transform -1 0 33120 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _442_
timestamp 1
transform -1 0 33764 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _443_
timestamp 1
transform 1 0 33120 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _444_
timestamp 1
transform 1 0 34132 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _445_
timestamp 1
transform 1 0 33580 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _446_
timestamp 1
transform 1 0 33396 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _447_
timestamp 1
transform 1 0 33120 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _448_
timestamp 1
transform 1 0 64768 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _449_
timestamp 1
transform 1 0 64768 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _450_
timestamp 1
transform -1 0 65412 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _451_
timestamp 1
transform 1 0 65320 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _452_
timestamp 1
transform -1 0 64676 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _453_
timestamp 1
transform 1 0 63848 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _454_
timestamp 1
transform -1 0 64676 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _455_
timestamp 1
transform 1 0 64676 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _456_
timestamp 1
transform -1 0 28888 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _457_
timestamp 1
transform 1 0 28060 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _458_
timestamp 1
transform 1 0 29900 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _459_
timestamp 1
transform 1 0 29532 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _460_
timestamp 1
transform 1 0 21712 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _461_
timestamp 1
transform 1 0 21528 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _462_
timestamp 1
transform 1 0 28980 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _463_
timestamp 1
transform 1 0 27508 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _464_
timestamp 1
transform -1 0 24840 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _465_
timestamp 1
transform 1 0 24288 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _466_
timestamp 1
transform -1 0 26312 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _467_
timestamp 1
transform 1 0 25668 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _468_
timestamp 1
transform 1 0 25668 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _469_
timestamp 1
transform 1 0 22908 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _470_
timestamp 1
transform 1 0 25208 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _471_
timestamp 1
transform 1 0 24656 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _472_
timestamp 1
transform 1 0 13524 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _473_
timestamp 1
transform 1 0 11776 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _474_
timestamp 1
transform 1 0 21804 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _475_
timestamp 1
transform -1 0 22080 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _476_
timestamp 1
transform 1 0 10948 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _477_
timestamp 1
transform 1 0 7912 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _478_
timestamp 1
transform 1 0 21252 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _479_
timestamp 1
transform 1 0 20884 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _480_
timestamp 1
transform -1 0 52072 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _481_
timestamp 1
transform 1 0 51244 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _482_
timestamp 1
transform 1 0 18124 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _483_
timestamp 1
transform -1 0 16008 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _484_
timestamp 1
transform 1 0 40112 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _485_
timestamp 1
transform 1 0 39100 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _486_
timestamp 1
transform 1 0 17388 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _487_
timestamp 1
transform 1 0 15180 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _488_
timestamp 1
transform 1 0 23828 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _489_
timestamp 1
transform 1 0 23092 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _490_
timestamp 1
transform 1 0 17572 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _491_
timestamp 1
transform 1 0 16468 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _492_
timestamp 1
transform 1 0 48392 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _493_
timestamp 1
transform -1 0 48668 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _494_
timestamp 1
transform 1 0 20056 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _495_
timestamp 1
transform 1 0 17756 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _496_
timestamp 1
transform 1 0 40112 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _497_
timestamp 1
transform 1 0 39284 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _498_
timestamp 1
transform -1 0 22816 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _499_
timestamp 1
transform 1 0 22080 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _500_
timestamp 1
transform 1 0 26404 0 -1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _501_
timestamp 1
transform 1 0 12144 0 -1 40800
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _502_
timestamp 1
transform 1 0 8372 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _503_
timestamp 1
transform 1 0 9476 0 1 39712
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _504_
timestamp 1
transform -1 0 22080 0 1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _505_
timestamp 1
transform 1 0 8740 0 -1 40800
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _506_
timestamp 1
transform -1 0 9200 0 -1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _507_
timestamp 1
transform 1 0 8464 0 1 38624
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _508_
timestamp 1
transform 1 0 7084 0 -1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _509_
timestamp 1
transform 1 0 8372 0 1 37536
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _510_
timestamp 1
transform 1 0 10580 0 1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _511_
timestamp 1
transform 1 0 10672 0 1 37536
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _512_
timestamp 1
transform 1 0 58512 0 -1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _513_
timestamp 1
transform -1 0 59892 0 -1 38624
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _514_
timestamp 1
transform 1 0 57868 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _515_
timestamp 1
transform 1 0 57592 0 -1 37536
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _516_
timestamp 1
transform 1 0 55016 0 1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _517_
timestamp 1
transform -1 0 57224 0 -1 38624
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _518_
timestamp 1
transform -1 0 54004 0 1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _519_
timestamp 1
transform -1 0 54648 0 1 37536
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _520_
timestamp 1
transform 1 0 54740 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _521_
timestamp 1
transform 1 0 54556 0 -1 40800
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _522_
timestamp 1
transform 1 0 52164 0 -1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _523_
timestamp 1
transform -1 0 54188 0 1 39712
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _524_
timestamp 1
transform 1 0 19044 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _525_
timestamp 1
transform 1 0 52164 0 -1 42976
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _526_
timestamp 1
transform 1 0 49588 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _527_
timestamp 1
transform 1 0 49404 0 -1 41888
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _528_
timestamp 1
transform 1 0 47656 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _529_
timestamp 1
transform -1 0 50600 0 -1 39712
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _530_
timestamp 1
transform 1 0 46460 0 1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _531_
timestamp 1
transform 1 0 46920 0 1 40800
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _532_
timestamp 1
transform 1 0 45080 0 -1 44064
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _533_
timestamp 1
transform 1 0 47012 0 1 42976
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _534_
timestamp 1
transform 1 0 44988 0 -1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _535_
timestamp 1
transform 1 0 45080 0 1 42976
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _536_
timestamp 1
transform 1 0 44804 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _537_
timestamp 1
transform 1 0 44804 0 -1 40800
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _538_
timestamp 1
transform 1 0 43792 0 -1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _539_
timestamp 1
transform -1 0 46368 0 1 37536
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _540_
timestamp 1
transform 1 0 41492 0 1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _541_
timestamp 1
transform -1 0 43792 0 -1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _542_
timestamp 1
transform 1 0 39744 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _543_
timestamp 1
transform -1 0 41768 0 -1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _544_
timestamp 1
transform -1 0 17388 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _545_
timestamp 1
transform 1 0 39284 0 1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _546_
timestamp 1
transform 1 0 37352 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _547_
timestamp 1
transform 1 0 39192 0 -1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _548_
timestamp 1
transform 1 0 34776 0 -1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _549_
timestamp 1
transform 1 0 35604 0 1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _550_
timestamp 1
transform 1 0 32016 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _551_
timestamp 1
transform -1 0 34960 0 -1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _552_
timestamp 1
transform 1 0 29716 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _553_
timestamp 1
transform 1 0 31556 0 -1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _554_
timestamp 1
transform 1 0 28888 0 -1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _555_
timestamp 1
transform 1 0 29900 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _556_
timestamp 1
transform 1 0 26772 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _557_
timestamp 1
transform 1 0 27600 0 -1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _558_
timestamp 1
transform 1 0 26496 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _559_
timestamp 1
transform 1 0 27048 0 -1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _560_
timestamp 1
transform 1 0 24104 0 -1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _561_
timestamp 1
transform 1 0 24656 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _562_
timestamp 1
transform 1 0 23460 0 -1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _563_
timestamp 1
transform 1 0 24564 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _564_
timestamp 1
transform -1 0 15548 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _565_
timestamp 1
transform 1 0 23828 0 1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _566_
timestamp 1
transform 1 0 19320 0 1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _567_
timestamp 1
transform 1 0 20608 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _568_
timestamp 1
transform 1 0 16652 0 -1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _569_
timestamp 1
transform 1 0 16744 0 -1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _570_
timestamp 1
transform 1 0 13524 0 -1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _571_
timestamp 1
transform 1 0 14904 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _572_
timestamp 1
transform -1 0 13800 0 -1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _573_
timestamp 1
transform 1 0 13524 0 1 38624
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _574_
timestamp 1
transform 1 0 9936 0 1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _575_
timestamp 1
transform 1 0 10672 0 1 42976
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _576_
timestamp 1
transform 1 0 12788 0 -1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _577_
timestamp 1
transform -1 0 15456 0 1 42976
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _578_
timestamp 1
transform 1 0 41860 0 -1 44064
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _579_
timestamp 1
transform -1 0 41308 0 -1 44064
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _580_
timestamp 1
transform 1 0 41860 0 -1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _581_
timestamp 1
transform 1 0 41676 0 1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _582_
timestamp 1
transform 1 0 42320 0 -1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _583_
timestamp 1
transform 1 0 42412 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _584_
timestamp 1
transform 1 0 15640 0 1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _585_
timestamp 1
transform -1 0 47932 0 1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _586_
timestamp 1
transform 1 0 50048 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _587_
timestamp 1
transform 1 0 49588 0 -1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _588_
timestamp 1
transform 1 0 63848 0 -1 35360
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _589_
timestamp 1
transform -1 0 64308 0 -1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _590_
timestamp 1
transform 1 0 64032 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _591_
timestamp 1
transform 1 0 64032 0 -1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _592_
timestamp 1
transform 1 0 64032 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _593_
timestamp 1
transform 1 0 64032 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _594_
timestamp 1
transform 1 0 64032 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _595_
timestamp 1
transform 1 0 64032 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _596_
timestamp 1
transform 1 0 64032 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _597_
timestamp 1
transform 1 0 64032 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _598_
timestamp 1
transform 1 0 64032 0 1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _599_
timestamp 1
transform 1 0 64032 0 1 23392
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _600_
timestamp 1
transform 1 0 64032 0 1 29920
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _601_
timestamp 1
transform 1 0 64032 0 1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _602_
timestamp 1
transform 1 0 63848 0 -1 36448
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _603_
timestamp 1
transform 1 0 64032 0 -1 33184
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _604_
timestamp 1
transform 1 0 18676 0 1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _605_
timestamp 1
transform 1 0 39928 0 -1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _606_
timestamp 1
transform 1 0 35052 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _607_
timestamp 1
transform 1 0 36708 0 -1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _608_
timestamp 1
transform -1 0 37812 0 1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _609_
timestamp 1
transform 1 0 34868 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _610_
timestamp 1
transform -1 0 38548 0 -1 44064
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _611_
timestamp 1
transform -1 0 38180 0 1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _612_
timestamp 1
transform 1 0 31648 0 -1 44064
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _613_
timestamp 1
transform 1 0 33488 0 -1 44064
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _614_
timestamp 1
transform -1 0 33212 0 1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _615_
timestamp 1
transform 1 0 31740 0 1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _616_
timestamp 1
transform 1 0 31740 0 -1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _617_
timestamp 1
transform -1 0 33396 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _618_
timestamp 1
transform 1 0 64032 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _619_
timestamp 1
transform 1 0 64032 0 1 12512
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _620_
timestamp 1
transform 1 0 63848 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _621_
timestamp 1
transform 1 0 63848 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _622_
timestamp 1
transform 1 0 27324 0 -1 44064
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _623_
timestamp 1
transform 1 0 29164 0 -1 44064
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _624_
timestamp 1
transform 1 0 20792 0 1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _625_
timestamp 1
transform 1 0 26588 0 1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _626_
timestamp 1
transform 1 0 23828 0 1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _627_
timestamp 1
transform 1 0 24012 0 -1 44064
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _628_
timestamp 1
transform 1 0 23000 0 -1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _629_
timestamp 1
transform 1 0 22816 0 -1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _630_
timestamp 1
transform 1 0 11500 0 -1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _631_
timestamp 1
transform 1 0 21712 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _632_
timestamp 1
transform 1 0 7728 0 -1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _633_
timestamp 1
transform -1 0 21068 0 -1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _634_
timestamp 1
transform 1 0 50600 0 1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _635_
timestamp 1
transform 1 0 16100 0 -1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _636_
timestamp 1
transform 1 0 38548 0 -1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _637_
timestamp 1
transform 1 0 14996 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _638_
timestamp 1
transform 1 0 21896 0 1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _639_
timestamp 1
transform 1 0 15364 0 1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _640_
timestamp 1
transform -1 0 48760 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _641_
timestamp 1
transform 1 0 17572 0 -1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _642_
timestamp 1
transform -1 0 40020 0 -1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _643_
timestamp 1
transform -1 0 21160 0 -1 44064
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  _666_
timestamp 1
transform 1 0 16100 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _667_
timestamp 1
transform -1 0 18584 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1
transform -1 0 64032 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1
transform -1 0 64768 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1
transform 1 0 64584 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1
transform 1 0 32936 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1
transform 1 0 34040 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1
transform 1 0 35788 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1
transform -1 0 37720 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1
transform 1 0 36708 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1
transform -1 0 37628 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1
transform -1 0 38364 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1
transform -1 0 20056 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1
transform 1 0 20056 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1
transform -1 0 64584 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1
transform -1 0 64676 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1
transform 1 0 64308 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1
transform -1 0 64768 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1
transform -1 0 64676 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1
transform -1 0 64860 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1
transform 1 0 64676 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1
transform -1 0 64676 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1
transform 1 0 49772 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1
transform -1 0 17572 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1
transform 1 0 17572 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1
transform -1 0 43240 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1
transform 1 0 43516 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1
transform -1 0 45448 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1
transform -1 0 17388 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1
transform -1 0 18124 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1
transform -1 0 25668 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1
transform -1 0 15180 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1
transform 1 0 45080 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1
transform 1 0 53820 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1
transform 1 0 53176 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ui_in[3]
timestamp 1
transform 1 0 35604 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ui_in[4]
timestamp 1
transform 1 0 36708 0 -1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_ui_in[3]
timestamp 1
transform 1 0 24656 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_ui_in[4]
timestamp 1
transform -1 0 28336 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_ui_in[3]
timestamp 1
transform 1 0 34776 0 -1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_ui_in[4]
timestamp 1
transform -1 0 38548 0 -1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_ui_in[3]
timestamp 1
transform -1 0 18584 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_ui_in[4]
timestamp 1
transform -1 0 18584 0 1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_ui_in[3]
timestamp 1
transform 1 0 19136 0 -1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_ui_in[4]
timestamp 1
transform -1 0 21712 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_ui_in[3]
timestamp 1
transform 1 0 63848 0 -1 31008
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_ui_in[4]
timestamp 1
transform 1 0 63848 0 1 31008
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_ui_in[3]
timestamp 1
transform 1 0 63848 0 -1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_ui_in[4]
timestamp 1
transform 1 0 63848 0 1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_ui_in[3]
timestamp 1
transform -1 0 43700 0 1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_ui_in[4]
timestamp 1
transform -1 0 42320 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_ui_in[3]
timestamp 1
transform 1 0 51428 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_ui_in[4]
timestamp 1
transform 1 0 50232 0 -1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinvlp_4  clkload0
timestamp 1
transform -1 0 26956 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkinvlp_4  clkload1
timestamp 1
transform 1 0 34500 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__bufinv_16  clkload2
timestamp 1
transform 1 0 17572 0 -1 38624
box -38 -48 2246 592
use sky130_fd_sc_hd__inv_6  clkload3
timestamp 1
transform 1 0 55568 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  clkload4
timestamp 1
transform 1 0 63848 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__clkinvlp_4  clkload5
timestamp 1
transform 1 0 51336 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__inv_4  clkload6
timestamp 1
transform 1 0 27140 0 -1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  clkload7
timestamp 1
transform 1 0 34868 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  clkload8
timestamp 1
transform 1 0 20148 0 -1 41888
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_4  clkload9
timestamp 1
transform -1 0 57776 0 -1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  clkload10
timestamp 1
transform -1 0 64308 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  clkload11
timestamp 1
transform 1 0 40480 0 -1 41888
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkload12
timestamp 1
transform 1 0 50692 0 1 39712
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout5
timestamp 1
transform -1 0 22632 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout6
timestamp 1
transform -1 0 35512 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout7
timestamp 1
transform 1 0 55660 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout8
timestamp 1
transform -1 0 57132 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout9
timestamp 1
transform -1 0 14168 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout10
timestamp 1
transform -1 0 15272 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout11
timestamp 1
transform 1 0 22632 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout12
timestamp 1
transform 1 0 27416 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout13
timestamp 1
transform -1 0 36248 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout14
timestamp 1
transform 1 0 35328 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout15
timestamp 1
transform -1 0 25576 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout16
timestamp 1
transform 1 0 63848 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout17
timestamp 1
transform -1 0 44252 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout18
timestamp 1
transform -1 0 41676 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout19
timestamp 1
transform -1 0 53544 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout20
timestamp 1
transform 1 0 53176 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout21
timestamp 1
transform 1 0 41860 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout22
timestamp 1
transform -1 0 23000 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout23
timestamp 1
transform -1 0 14720 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout24
timestamp 1
transform -1 0 21712 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout25
timestamp 1
transform -1 0 13432 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout26
timestamp 1
transform 1 0 28980 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout27
timestamp 1
transform 1 0 31188 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout28
timestamp 1
transform 1 0 33580 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout29
timestamp 1
transform -1 0 26312 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout30
timestamp 1
transform 1 0 64860 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout31
timestamp 1
transform 1 0 41216 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout32
timestamp 1
transform -1 0 41216 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout33
timestamp 1
transform -1 0 41676 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout34
timestamp 1
transform -1 0 52716 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout35
timestamp 1
transform 1 0 53728 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout36
timestamp 1
transform 1 0 44436 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout37
timestamp 1
transform -1 0 12512 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout38
timestamp 1
transform -1 0 13616 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout39
timestamp 1
transform -1 0 13248 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout40
timestamp 1
transform -1 0 19228 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout41
timestamp 1
transform -1 0 23368 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 1
transform -1 0 29532 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout43
timestamp 1
transform -1 0 32660 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout44
timestamp 1
transform 1 0 30360 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout45
timestamp 1
transform -1 0 31924 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout46
timestamp 1
transform 1 0 65228 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout47
timestamp 1
transform -1 0 39836 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout48
timestamp 1
transform -1 0 44620 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout49
timestamp 1
transform 1 0 39284 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout50
timestamp 1
transform -1 0 47564 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout51
timestamp 1
transform -1 0 46920 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout52
timestamp 1
transform 1 0 53544 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout53
timestamp 1
transform -1 0 54096 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout54
timestamp 1
transform 1 0 52716 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout55
timestamp 1
transform 1 0 38548 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout56
timestamp 1
transform 1 0 31924 0 1 44064
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_688
timestamp 1636968456
transform 1 0 63848 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_700
timestamp 1
transform 1 0 64952 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_704
timestamp 1
transform 1 0 65320 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_688
timestamp 1
transform 1 0 63848 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_707
timestamp 1
transform 1 0 65596 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_688
timestamp 1
transform 1 0 63848 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_707
timestamp 1
transform 1 0 65596 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_4_710
timestamp 1
transform 1 0 65872 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_706
timestamp 1
transform 1 0 65504 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_712
timestamp 1
transform 1 0 66056 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_708
timestamp 1
transform 1 0 65688 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_712
timestamp 1
transform 1 0 66056 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_708
timestamp 1
transform 1 0 65688 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_712
timestamp 1
transform 1 0 66056 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_688
timestamp 1
transform 1 0 63848 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_710
timestamp 1
transform 1 0 65872 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_699
timestamp 1636968456
transform 1 0 64860 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_711
timestamp 1
transform 1 0 65964 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_706
timestamp 1
transform 1 0 65504 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_712
timestamp 1
transform 1 0 66056 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_694
timestamp 1
transform 1 0 64400 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_708
timestamp 1
transform 1 0 65688 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_712
timestamp 1
transform 1 0 66056 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_688
timestamp 1
transform 1 0 63848 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_694
timestamp 1
transform 1 0 64400 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_704
timestamp 1
transform 1 0 65320 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_688
timestamp 1
transform 1 0 63848 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_710
timestamp 1
transform 1 0 65872 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_688
timestamp 1
transform 1 0 63848 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_688
timestamp 1
transform 1 0 63848 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_705
timestamp 1
transform 1 0 65412 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_688
timestamp 1
transform 1 0 63848 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_688
timestamp 1
transform 1 0 63848 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_710
timestamp 1
transform 1 0 65872 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_688
timestamp 1
transform 1 0 63848 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_705
timestamp 1
transform 1 0 65412 0 1 10336
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_688
timestamp 1636968456
transform 1 0 63848 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_700
timestamp 1
transform 1 0 64952 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_704
timestamp 1
transform 1 0 65320 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_688
timestamp 1
transform 1 0 63848 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_694
timestamp 1
transform 1 0 64400 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_688
timestamp 1
transform 1 0 63848 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_710
timestamp 1
transform 1 0 65872 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_688
timestamp 1
transform 1 0 63848 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_688
timestamp 1636968456
transform 1 0 63848 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_700
timestamp 1636968456
transform 1 0 64952 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_712
timestamp 1
transform 1 0 66056 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_688
timestamp 1636968456
transform 1 0 63848 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_700
timestamp 1636968456
transform 1 0 64952 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_712
timestamp 1
transform 1 0 66056 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_688
timestamp 1636968456
transform 1 0 63848 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_700
timestamp 1636968456
transform 1 0 64952 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_712
timestamp 1
transform 1 0 66056 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_688
timestamp 1
transform 1 0 63848 0 1 14688
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_698
timestamp 1636968456
transform 1 0 64768 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_710
timestamp 1
transform 1 0 65872 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_688
timestamp 1
transform 1 0 63848 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_705
timestamp 1
transform 1 0 65412 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_688
timestamp 1
transform 1 0 63848 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_710
timestamp 1
transform 1 0 65872 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_688
timestamp 1
transform 1 0 63848 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_688
timestamp 1
transform 1 0 63848 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_694
timestamp 1
transform 1 0 64400 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_697
timestamp 1636968456
transform 1 0 64676 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_709
timestamp 1
transform 1 0 65780 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_688
timestamp 1
transform 1 0 63848 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_694
timestamp 1
transform 1 0 64400 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_688
timestamp 1
transform 1 0 63848 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_710
timestamp 1
transform 1 0 65872 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_688
timestamp 1
transform 1 0 63848 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_688
timestamp 1
transform 1 0 63848 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_688
timestamp 1
transform 1 0 63848 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_710
timestamp 1
transform 1 0 65872 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_688
timestamp 1
transform 1 0 63848 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_705
timestamp 1
transform 1 0 65412 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_688
timestamp 1
transform 1 0 63848 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_705
timestamp 1
transform 1 0 65412 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_688
timestamp 1
transform 1 0 63848 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_696
timestamp 1
transform 1 0 64584 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_688
timestamp 1
transform 1 0 63848 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_710
timestamp 1
transform 1 0 65872 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_697
timestamp 1
transform 1 0 64676 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_709
timestamp 1
transform 1 0 65780 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_688
timestamp 1
transform 1 0 63848 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_692
timestamp 1
transform 1 0 64216 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_704
timestamp 1
transform 1 0 65320 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_712
timestamp 1
transform 1 0 66056 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_688
timestamp 1
transform 1 0 63848 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_710
timestamp 1
transform 1 0 65872 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_708
timestamp 1
transform 1 0 65688 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_712
timestamp 1
transform 1 0 66056 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_708
timestamp 1
transform 1 0 65688 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_712
timestamp 1
transform 1 0 66056 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_693
timestamp 1
transform 1 0 64308 0 -1 25568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_688
timestamp 1636968456
transform 1 0 63848 0 1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_700
timestamp 1636968456
transform 1 0 64952 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_712
timestamp 1
transform 1 0 66056 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_688
timestamp 1
transform 1 0 63848 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_688
timestamp 1
transform 1 0 63848 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_710
timestamp 1
transform 1 0 65872 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_688
timestamp 1
transform 1 0 63848 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_705
timestamp 1
transform 1 0 65412 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_50_688
timestamp 1
transform 1 0 63848 0 1 27744
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_696
timestamp 1636968456
transform 1 0 64584 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_708
timestamp 1
transform 1 0 65688 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_712
timestamp 1
transform 1 0 66056 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_688
timestamp 1
transform 1 0 63848 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_703
timestamp 1
transform 1 0 65228 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_688
timestamp 1
transform 1 0 63848 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_710
timestamp 1
transform 1 0 65872 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_688
timestamp 1
transform 1 0 63848 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_694
timestamp 1
transform 1 0 64400 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_688
timestamp 1
transform 1 0 63848 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_710
timestamp 1
transform 1 0 65872 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_708
timestamp 1
transform 1 0 65688 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_712
timestamp 1
transform 1 0 66056 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_708
timestamp 1
transform 1 0 65688 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_712
timestamp 1
transform 1 0 66056 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_688
timestamp 1
transform 1 0 63848 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_688
timestamp 1
transform 1 0 63848 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_692
timestamp 1
transform 1 0 64216 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_702
timestamp 1
transform 1 0 65136 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_710
timestamp 1
transform 1 0 65872 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_688
timestamp 1
transform 1 0 63848 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_710
timestamp 1
transform 1 0 65872 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_688
timestamp 1
transform 1 0 63848 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_694
timestamp 1
transform 1 0 64400 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_704
timestamp 1
transform 1 0 65320 0 1 33184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_688
timestamp 1636968456
transform 1 0 63848 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_700
timestamp 1
transform 1 0 64952 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_710
timestamp 1
transform 1 0 65872 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_706
timestamp 1
transform 1 0 65504 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_712
timestamp 1
transform 1 0 66056 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_708
timestamp 1
transform 1 0 65688 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_712
timestamp 1
transform 1 0 66056 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_688
timestamp 1
transform 1 0 63848 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_710
timestamp 1
transform 1 0 65872 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_708
timestamp 1
transform 1 0 65688 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_712
timestamp 1
transform 1 0 66056 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_706
timestamp 1
transform 1 0 65504 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_712
timestamp 1
transform 1 0 66056 0 1 36448
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1636968456
transform 1 0 828 0 -1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1636968456
transform 1 0 1932 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_27
timestamp 1
transform 1 0 3036 0 -1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_29
timestamp 1636968456
transform 1 0 3220 0 -1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_41
timestamp 1636968456
transform 1 0 4324 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_53
timestamp 1
transform 1 0 5428 0 -1 37536
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1636968456
transform 1 0 5796 0 -1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1636968456
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_81
timestamp 1
transform 1 0 8004 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_67_85
timestamp 1
transform 1 0 8372 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_91
timestamp 1
transform 1 0 8924 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_101
timestamp 1
transform 1 0 9844 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_109
timestamp 1
transform 1 0 10580 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_122
timestamp 1
transform 1 0 11776 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_126
timestamp 1
transform 1 0 12144 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_136
timestamp 1
transform 1 0 13064 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1
transform 1 0 15364 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1
transform 1 0 15916 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_169
timestamp 1
transform 1 0 16100 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_175
timestamp 1
transform 1 0 16652 0 -1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_206
timestamp 1636968456
transform 1 0 19504 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_218
timestamp 1
transform 1 0 20608 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_225
timestamp 1
transform 1 0 21252 0 -1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_235
timestamp 1636968456
transform 1 0 22172 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_247
timestamp 1
transform 1 0 23276 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_251
timestamp 1
transform 1 0 23644 0 -1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_253
timestamp 1636968456
transform 1 0 23828 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_265
timestamp 1
transform 1 0 24932 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_67_290
timestamp 1
transform 1 0 27232 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_296
timestamp 1
transform 1 0 27784 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_306
timestamp 1
transform 1 0 28704 0 -1 37536
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_309
timestamp 1636968456
transform 1 0 28980 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_321
timestamp 1
transform 1 0 30084 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_333
timestamp 1
transform 1 0 31188 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_67_345
timestamp 1
transform 1 0 32292 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_365
timestamp 1
transform 1 0 34132 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_371
timestamp 1
transform 1 0 34684 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_413
timestamp 1
transform 1 0 38548 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_419
timestamp 1
transform 1 0 39100 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_421
timestamp 1
transform 1 0 39284 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_427
timestamp 1
transform 1 0 39836 0 -1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1636968456
transform 1 0 41860 0 -1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1636968456
transform 1 0 42964 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_473
timestamp 1
transform 1 0 44068 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_495
timestamp 1
transform 1 0 46092 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1
transform 1 0 46828 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_523
timestamp 1
transform 1 0 48668 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_531
timestamp 1
transform 1 0 49404 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_533
timestamp 1
transform 1 0 49588 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_546
timestamp 1
transform 1 0 50784 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_556
timestamp 1
transform 1 0 51704 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_570
timestamp 1
transform 1 0 52992 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_583
timestamp 1
transform 1 0 54188 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_587
timestamp 1
transform 1 0 54556 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_589
timestamp 1
transform 1 0 54740 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_597
timestamp 1
transform 1 0 55476 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_605
timestamp 1
transform 1 0 56212 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_67_617
timestamp 1
transform 1 0 57316 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_67_643
timestamp 1
transform 1 0 59708 0 -1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_645
timestamp 1636968456
transform 1 0 59892 0 -1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_657
timestamp 1636968456
transform 1 0 60996 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_669
timestamp 1
transform 1 0 62100 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_67_693
timestamp 1
transform 1 0 64308 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_699
timestamp 1
transform 1 0 64860 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_701
timestamp 1
transform 1 0 65044 0 -1 37536
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1636968456
transform 1 0 828 0 1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1636968456
transform 1 0 1932 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1
transform 1 0 3036 0 1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1636968456
transform 1 0 3220 0 1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1636968456
transform 1 0 4324 0 1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1636968456
transform 1 0 5428 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_65
timestamp 1
transform 1 0 6532 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_73
timestamp 1
transform 1 0 7268 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_108
timestamp 1
transform 1 0 10488 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1
transform 1 0 12788 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1
transform 1 0 13340 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_141
timestamp 1
transform 1 0 13524 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_68_206
timestamp 1
transform 1 0 19504 0 1 37536
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_238
timestamp 1636968456
transform 1 0 22448 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_250
timestamp 1
transform 1 0 23552 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_302
timestamp 1
transform 1 0 28336 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_68_317
timestamp 1
transform 1 0 29716 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_68_339
timestamp 1
transform 1 0 31740 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_362
timestamp 1
transform 1 0 33856 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_380
timestamp 1
transform 1 0 35512 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_401
timestamp 1
transform 1 0 37444 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_439
timestamp 1
transform 1 0 40940 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_68_450
timestamp 1
transform 1 0 41952 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1
transform 1 0 43700 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1
transform 1 0 44252 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_498
timestamp 1
transform 1 0 46368 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_533
timestamp 1
transform 1 0 49588 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_537
timestamp 1
transform 1 0 49956 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_558
timestamp 1
transform 1 0 51888 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_564
timestamp 1
transform 1 0 52440 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_589
timestamp 1
transform 1 0 54740 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_613
timestamp 1
transform 1 0 56948 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_643
timestamp 1
transform 1 0 59708 0 1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_654
timestamp 1636968456
transform 1 0 60720 0 1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_666
timestamp 1636968456
transform 1 0 61824 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_678
timestamp 1
transform 1 0 62928 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_682
timestamp 1
transform 1 0 63296 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_691
timestamp 1
transform 1 0 64124 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_699
timestamp 1
transform 1 0 64860 0 1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_701
timestamp 1636968456
transform 1 0 65044 0 1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1636968456
transform 1 0 828 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1636968456
transform 1 0 1932 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1636968456
transform 1 0 3036 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1636968456
transform 1 0 4140 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1
transform 1 0 5244 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1
transform 1 0 5612 0 -1 38624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1636968456
transform 1 0 5796 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_69
timestamp 1
transform 1 0 6900 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_69_91
timestamp 1
transform 1 0 8924 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_113
timestamp 1
transform 1 0 10948 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_132
timestamp 1
transform 1 0 12696 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_140
timestamp 1
transform 1 0 13432 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_69_152
timestamp 1
transform 1 0 14536 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_158
timestamp 1
transform 1 0 15088 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_178
timestamp 1
transform 1 0 16928 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_184
timestamp 1
transform 1 0 17480 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_218
timestamp 1
transform 1 0 20608 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_240
timestamp 1
transform 1 0 22632 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_244
timestamp 1
transform 1 0 23000 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_254
timestamp 1
transform 1 0 23920 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_276
timestamp 1
transform 1 0 25944 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_281
timestamp 1
transform 1 0 26404 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_287
timestamp 1
transform 1 0 26956 0 -1 38624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1636968456
transform 1 0 31556 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_349
timestamp 1
transform 1 0 32660 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_353
timestamp 1
transform 1 0 33028 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_402
timestamp 1
transform 1 0 37536 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_408
timestamp 1
transform 1 0 38088 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_429
timestamp 1
transform 1 0 40020 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_442
timestamp 1
transform 1 0 41216 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_449
timestamp 1
transform 1 0 41860 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_498
timestamp 1
transform 1 0 46368 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_69_514
timestamp 1
transform 1 0 47840 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_529
timestamp 1
transform 1 0 49220 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1
transform 1 0 51428 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1
transform 1 0 51980 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_578
timestamp 1
transform 1 0 53728 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_590
timestamp 1
transform 1 0 54832 0 -1 38624
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_654
timestamp 1636968456
transform 1 0 60720 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_666
timestamp 1
transform 1 0 61824 0 -1 38624
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_673
timestamp 1636968456
transform 1 0 62468 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_685
timestamp 1636968456
transform 1 0 63572 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_697
timestamp 1636968456
transform 1 0 64676 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_709
timestamp 1
transform 1 0 65780 0 -1 38624
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1636968456
transform 1 0 828 0 1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1636968456
transform 1 0 1932 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1
transform 1 0 3036 0 1 38624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1636968456
transform 1 0 3220 0 1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1636968456
transform 1 0 4324 0 1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1636968456
transform 1 0 5428 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_65
timestamp 1
transform 1 0 6532 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_73
timestamp 1
transform 1 0 7268 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_70_85
timestamp 1
transform 1 0 8372 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_129
timestamp 1
transform 1 0 12420 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_170
timestamp 1
transform 1 0 16192 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_70_197
timestamp 1
transform 1 0 18676 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_203
timestamp 1
transform 1 0 19228 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_282
timestamp 1
transform 1 0 26496 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_70_306
timestamp 1
transform 1 0 28704 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_309
timestamp 1
transform 1 0 28980 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_333
timestamp 1
transform 1 0 31188 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_354
timestamp 1
transform 1 0 33120 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_439
timestamp 1
transform 1 0 40940 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_70_473
timestamp 1
transform 1 0 44068 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_70_494
timestamp 1
transform 1 0 46000 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_515
timestamp 1
transform 1 0 47932 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_533
timestamp 1
transform 1 0 49588 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_70_545
timestamp 1
transform 1 0 50692 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_555
timestamp 1
transform 1 0 51612 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1
transform 1 0 54004 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1
transform 1 0 54556 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_589
timestamp 1
transform 1 0 54740 0 1 38624
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_612
timestamp 1636968456
transform 1 0 56856 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_624
timestamp 1
transform 1 0 57960 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_643
timestamp 1
transform 1 0 59708 0 1 38624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_653
timestamp 1636968456
transform 1 0 60628 0 1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_665
timestamp 1636968456
transform 1 0 61732 0 1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_677
timestamp 1636968456
transform 1 0 62836 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_689
timestamp 1
transform 1 0 63940 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_697
timestamp 1
transform 1 0 64676 0 1 38624
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_701
timestamp 1636968456
transform 1 0 65044 0 1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1636968456
transform 1 0 828 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1636968456
transform 1 0 1932 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1636968456
transform 1 0 3036 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1636968456
transform 1 0 4140 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1
transform 1 0 5244 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1
transform 1 0 5612 0 -1 39712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1636968456
transform 1 0 5796 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_69
timestamp 1
transform 1 0 6900 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_73
timestamp 1
transform 1 0 7268 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_103
timestamp 1
transform 1 0 10028 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1
transform 1 0 10764 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_122
timestamp 1
transform 1 0 11776 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_153
timestamp 1
transform 1 0 14628 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_71_169
timestamp 1
transform 1 0 16100 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_71_195
timestamp 1
transform 1 0 18492 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_201
timestamp 1
transform 1 0 19044 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_222
timestamp 1
transform 1 0 20976 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_243
timestamp 1
transform 1 0 22908 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_71_260
timestamp 1
transform 1 0 24472 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_266
timestamp 1
transform 1 0 25024 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_276
timestamp 1
transform 1 0 25944 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_297
timestamp 1
transform 1 0 27876 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_71_320
timestamp 1
transform 1 0 29992 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_326
timestamp 1
transform 1 0 30544 0 -1 39712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_366
timestamp 1636968456
transform 1 0 34224 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_378
timestamp 1
transform 1 0 35328 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_382
timestamp 1
transform 1 0 35696 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_422
timestamp 1
transform 1 0 39376 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_71_449
timestamp 1
transform 1 0 41860 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_478
timestamp 1
transform 1 0 44528 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_71_513
timestamp 1
transform 1 0 47748 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_558
timestamp 1
transform 1 0 51888 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_561
timestamp 1
transform 1 0 52164 0 -1 39712
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_580
timestamp 1636968456
transform 1 0 53912 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_592
timestamp 1
transform 1 0 55016 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_596
timestamp 1
transform 1 0 55384 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_606
timestamp 1
transform 1 0 56304 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1
transform 1 0 57132 0 -1 39712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_617
timestamp 1636968456
transform 1 0 57316 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_629
timestamp 1
transform 1 0 58420 0 -1 39712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_658
timestamp 1636968456
transform 1 0 61088 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_670
timestamp 1
transform 1 0 62192 0 -1 39712
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_673
timestamp 1636968456
transform 1 0 62468 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_685
timestamp 1636968456
transform 1 0 63572 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_697
timestamp 1636968456
transform 1 0 64676 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_709
timestamp 1
transform 1 0 65780 0 -1 39712
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1636968456
transform 1 0 828 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1636968456
transform 1 0 1932 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1
transform 1 0 3036 0 1 39712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1636968456
transform 1 0 3220 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1636968456
transform 1 0 4324 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1636968456
transform 1 0 5428 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_65
timestamp 1
transform 1 0 6532 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_73
timestamp 1
transform 1 0 7268 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_85
timestamp 1
transform 1 0 8372 0 1 39712
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_120
timestamp 1636968456
transform 1 0 11592 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_141
timestamp 1
transform 1 0 13524 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_183
timestamp 1
transform 1 0 17388 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_194
timestamp 1
transform 1 0 18400 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_197
timestamp 1
transform 1 0 18676 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_230
timestamp 1
transform 1 0 21712 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_248
timestamp 1
transform 1 0 23368 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_281
timestamp 1
transform 1 0 26404 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_72_305
timestamp 1
transform 1 0 28612 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_72_309
timestamp 1
transform 1 0 28980 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1
transform 1 0 33396 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1
transform 1 0 33948 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_374
timestamp 1
transform 1 0 34960 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_395
timestamp 1
transform 1 0 36892 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_399
timestamp 1
transform 1 0 37260 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_421
timestamp 1
transform 1 0 39284 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_425
timestamp 1
transform 1 0 39652 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_455
timestamp 1
transform 1 0 42412 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_461
timestamp 1
transform 1 0 42964 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_72_473
timestamp 1
transform 1 0 44068 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_477
timestamp 1
transform 1 0 44436 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_72_509
timestamp 1
transform 1 0 47380 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_542
timestamp 1
transform 1 0 50416 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_556
timestamp 1
transform 1 0 51704 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_583
timestamp 1
transform 1 0 54188 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1
transform 1 0 54556 0 1 39712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_607
timestamp 1636968456
transform 1 0 56396 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_619
timestamp 1636968456
transform 1 0 57500 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_631
timestamp 1636968456
transform 1 0 58604 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_643
timestamp 1
transform 1 0 59708 0 1 39712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_645
timestamp 1636968456
transform 1 0 59892 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_657
timestamp 1636968456
transform 1 0 60996 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_669
timestamp 1636968456
transform 1 0 62100 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_681
timestamp 1636968456
transform 1 0 63204 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_693
timestamp 1
transform 1 0 64308 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_699
timestamp 1
transform 1 0 64860 0 1 39712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_701
timestamp 1636968456
transform 1 0 65044 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1636968456
transform 1 0 828 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1636968456
transform 1 0 1932 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1636968456
transform 1 0 3036 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1636968456
transform 1 0 4140 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1
transform 1 0 5244 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1
transform 1 0 5612 0 -1 40800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1636968456
transform 1 0 5796 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_69
timestamp 1
transform 1 0 6900 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_77
timestamp 1
transform 1 0 7636 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_122
timestamp 1
transform 1 0 11776 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_149
timestamp 1
transform 1 0 14260 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_73_200
timestamp 1
transform 1 0 18952 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1
transform 1 0 21068 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_248
timestamp 1
transform 1 0 23368 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_278
timestamp 1
transform 1 0 26128 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_323
timestamp 1
transform 1 0 30268 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_337
timestamp 1
transform 1 0 31556 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_368
timestamp 1
transform 1 0 34408 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_413
timestamp 1
transform 1 0 38548 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_419
timestamp 1
transform 1 0 39100 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_453
timestamp 1
transform 1 0 42228 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_474
timestamp 1
transform 1 0 44160 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_480
timestamp 1
transform 1 0 44712 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_502
timestamp 1
transform 1 0 46736 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_505
timestamp 1
transform 1 0 47012 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_518
timestamp 1
transform 1 0 48208 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_581
timestamp 1
transform 1 0 54004 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_73_610
timestamp 1
transform 1 0 56672 0 -1 40800
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_617
timestamp 1636968456
transform 1 0 57316 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_629
timestamp 1636968456
transform 1 0 58420 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_641
timestamp 1636968456
transform 1 0 59524 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_653
timestamp 1636968456
transform 1 0 60628 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_665
timestamp 1
transform 1 0 61732 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_671
timestamp 1
transform 1 0 62284 0 -1 40800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_673
timestamp 1636968456
transform 1 0 62468 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_685
timestamp 1636968456
transform 1 0 63572 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_697
timestamp 1636968456
transform 1 0 64676 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_709
timestamp 1
transform 1 0 65780 0 -1 40800
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1636968456
transform 1 0 828 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1636968456
transform 1 0 1932 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1
transform 1 0 3036 0 1 40800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1636968456
transform 1 0 3220 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1636968456
transform 1 0 4324 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1636968456
transform 1 0 5428 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_65
timestamp 1
transform 1 0 6532 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_73
timestamp 1
transform 1 0 7268 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_114
timestamp 1
transform 1 0 11040 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_74_150
timestamp 1
transform 1 0 14352 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_156
timestamp 1
transform 1 0 14904 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_177
timestamp 1
transform 1 0 16836 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_192
timestamp 1
transform 1 0 18216 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_206
timestamp 1
transform 1 0 19504 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_250
timestamp 1
transform 1 0 23552 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_302
timestamp 1
transform 1 0 28336 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_74_326
timestamp 1
transform 1 0 30544 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_342
timestamp 1
transform 1 0 32016 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1
transform 1 0 33948 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_395
timestamp 1
transform 1 0 36892 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_74_417
timestamp 1
transform 1 0 38916 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_430
timestamp 1
transform 1 0 40112 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_454
timestamp 1
transform 1 0 42320 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1
transform 1 0 44252 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_486
timestamp 1
transform 1 0 45264 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1
transform 1 0 48852 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1
transform 1 0 49404 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_582
timestamp 1
transform 1 0 54096 0 1 40800
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_620
timestamp 1636968456
transform 1 0 57592 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_632
timestamp 1636968456
transform 1 0 58696 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_645
timestamp 1636968456
transform 1 0 59892 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_657
timestamp 1636968456
transform 1 0 60996 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_669
timestamp 1636968456
transform 1 0 62100 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_681
timestamp 1636968456
transform 1 0 63204 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_693
timestamp 1
transform 1 0 64308 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_699
timestamp 1
transform 1 0 64860 0 1 40800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_701
timestamp 1636968456
transform 1 0 65044 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1636968456
transform 1 0 828 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1636968456
transform 1 0 1932 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1636968456
transform 1 0 3036 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1636968456
transform 1 0 4140 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1
transform 1 0 5244 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1
transform 1 0 5612 0 -1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1636968456
transform 1 0 5796 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_69
timestamp 1
transform 1 0 6900 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_77
timestamp 1
transform 1 0 7636 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_107
timestamp 1
transform 1 0 10396 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1
transform 1 0 10764 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_113
timestamp 1
transform 1 0 10948 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_147
timestamp 1
transform 1 0 14076 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_169
timestamp 1
transform 1 0 16100 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_175
timestamp 1
transform 1 0 16652 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_204
timestamp 1
transform 1 0 19320 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_243
timestamp 1
transform 1 0 22908 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_264
timestamp 1
transform 1 0 24840 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_75_277
timestamp 1
transform 1 0 26036 0 -1 41888
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_318
timestamp 1636968456
transform 1 0 29808 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_330
timestamp 1
transform 1 0 30912 0 -1 41888
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1636968456
transform 1 0 31556 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_349
timestamp 1
transform 1 0 32660 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_75_361
timestamp 1
transform 1 0 33764 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_75_366
timestamp 1
transform 1 0 34224 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_75_404
timestamp 1
transform 1 0 37720 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_433
timestamp 1
transform 1 0 40388 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_75_445
timestamp 1
transform 1 0 41492 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_486
timestamp 1
transform 1 0 45264 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_490
timestamp 1
transform 1 0 45632 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_500
timestamp 1
transform 1 0 46552 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_75_505
timestamp 1
transform 1 0 47012 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_526
timestamp 1
transform 1 0 48944 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_530
timestamp 1
transform 1 0 49312 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_554
timestamp 1
transform 1 0 51520 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_586
timestamp 1
transform 1 0 54464 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_75_599
timestamp 1
transform 1 0 55660 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_75_610
timestamp 1
transform 1 0 56672 0 -1 41888
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_617
timestamp 1636968456
transform 1 0 57316 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_629
timestamp 1636968456
transform 1 0 58420 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_641
timestamp 1636968456
transform 1 0 59524 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_653
timestamp 1636968456
transform 1 0 60628 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_665
timestamp 1
transform 1 0 61732 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_671
timestamp 1
transform 1 0 62284 0 -1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_673
timestamp 1636968456
transform 1 0 62468 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_685
timestamp 1636968456
transform 1 0 63572 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_697
timestamp 1636968456
transform 1 0 64676 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_709
timestamp 1
transform 1 0 65780 0 -1 41888
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1636968456
transform 1 0 828 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1636968456
transform 1 0 1932 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1
transform 1 0 3036 0 1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1636968456
transform 1 0 3220 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1636968456
transform 1 0 4324 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1636968456
transform 1 0 5428 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1636968456
transform 1 0 6532 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1
transform 1 0 7636 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1
transform 1 0 8188 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_85
timestamp 1
transform 1 0 8372 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_91
timestamp 1
transform 1 0 8924 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_100
timestamp 1
transform 1 0 9752 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_122
timestamp 1
transform 1 0 11776 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1
transform 1 0 13340 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_141
timestamp 1
transform 1 0 13524 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_159
timestamp 1
transform 1 0 15180 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_181
timestamp 1
transform 1 0 17204 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_194
timestamp 1
transform 1 0 18400 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_197
timestamp 1
transform 1 0 18676 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_210
timestamp 1
transform 1 0 19872 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_253
timestamp 1
transform 1 0 23828 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_76_264
timestamp 1
transform 1 0 24840 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_270
timestamp 1
transform 1 0 25392 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_282
timestamp 1
transform 1 0 26496 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_303
timestamp 1
transform 1 0 28428 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1
transform 1 0 28796 0 1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_315
timestamp 1636968456
transform 1 0 29532 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_327
timestamp 1
transform 1 0 30636 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_76_377
timestamp 1
transform 1 0 35236 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_76_414
timestamp 1
transform 1 0 38640 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_76_447
timestamp 1
transform 1 0 41676 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1
transform 1 0 43700 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1
transform 1 0 44252 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_488
timestamp 1
transform 1 0 45448 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_498
timestamp 1
transform 1 0 46368 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_519
timestamp 1
transform 1 0 48300 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_528
timestamp 1
transform 1 0 49128 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_569
timestamp 1
transform 1 0 52900 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_582
timestamp 1
transform 1 0 54096 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_76_589
timestamp 1
transform 1 0 54740 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_597
timestamp 1
transform 1 0 55476 0 1 41888
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_605
timestamp 1636968456
transform 1 0 56212 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_617
timestamp 1636968456
transform 1 0 57316 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_629
timestamp 1636968456
transform 1 0 58420 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_641
timestamp 1
transform 1 0 59524 0 1 41888
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_645
timestamp 1636968456
transform 1 0 59892 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_657
timestamp 1636968456
transform 1 0 60996 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_669
timestamp 1636968456
transform 1 0 62100 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_681
timestamp 1636968456
transform 1 0 63204 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_693
timestamp 1
transform 1 0 64308 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_699
timestamp 1
transform 1 0 64860 0 1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_701
timestamp 1636968456
transform 1 0 65044 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1636968456
transform 1 0 828 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1636968456
transform 1 0 1932 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1636968456
transform 1 0 3036 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1636968456
transform 1 0 4140 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1
transform 1 0 5244 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1
transform 1 0 5612 0 -1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1636968456
transform 1 0 5796 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1636968456
transform 1 0 6900 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_81
timestamp 1
transform 1 0 8004 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_89
timestamp 1
transform 1 0 8740 0 -1 42976
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_99
timestamp 1636968456
transform 1 0 9660 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1
transform 1 0 10764 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_113
timestamp 1
transform 1 0 10948 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_126
timestamp 1
transform 1 0 12144 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_132
timestamp 1
transform 1 0 12696 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_153
timestamp 1
transform 1 0 14628 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_205
timestamp 1
transform 1 0 19412 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_209
timestamp 1
transform 1 0 19780 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_77_221
timestamp 1
transform 1 0 20884 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_77_318
timestamp 1
transform 1 0 29808 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_328
timestamp 1
transform 1 0 30728 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_363
timestamp 1
transform 1 0 33948 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_373
timestamp 1
transform 1 0 34868 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_381
timestamp 1
transform 1 0 35604 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_418
timestamp 1
transform 1 0 39008 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_428
timestamp 1
transform 1 0 39928 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_478
timestamp 1
transform 1 0 44528 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_482
timestamp 1
transform 1 0 44896 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1
transform 1 0 46828 0 -1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_531
timestamp 1636968456
transform 1 0 49404 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_543
timestamp 1
transform 1 0 50508 0 -1 42976
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_77_584
timestamp 1636968456
transform 1 0 54280 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_596
timestamp 1636968456
transform 1 0 55384 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_608
timestamp 1
transform 1 0 56488 0 -1 42976
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_77_617
timestamp 1636968456
transform 1 0 57316 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_629
timestamp 1636968456
transform 1 0 58420 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_641
timestamp 1636968456
transform 1 0 59524 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_653
timestamp 1636968456
transform 1 0 60628 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_665
timestamp 1
transform 1 0 61732 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_671
timestamp 1
transform 1 0 62284 0 -1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_673
timestamp 1636968456
transform 1 0 62468 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_685
timestamp 1636968456
transform 1 0 63572 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_697
timestamp 1636968456
transform 1 0 64676 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_709
timestamp 1
transform 1 0 65780 0 -1 42976
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1636968456
transform 1 0 828 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1636968456
transform 1 0 1932 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1
transform 1 0 3036 0 1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1636968456
transform 1 0 3220 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1636968456
transform 1 0 4324 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1636968456
transform 1 0 5428 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1636968456
transform 1 0 6532 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1
transform 1 0 7636 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1
transform 1 0 8188 0 1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1636968456
transform 1 0 8372 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1636968456
transform 1 0 9476 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_109
timestamp 1
transform 1 0 10580 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_131
timestamp 1
transform 1 0 12604 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1
transform 1 0 13340 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_162
timestamp 1
transform 1 0 15456 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_78_217
timestamp 1
transform 1 0 20516 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_78_282
timestamp 1
transform 1 0 26496 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_298
timestamp 1
transform 1 0 27968 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_78_330
timestamp 1
transform 1 0 30912 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1
transform 1 0 33948 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_383
timestamp 1
transform 1 0 35788 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_78_418
timestamp 1
transform 1 0 39008 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_78_425
timestamp 1
transform 1 0 39652 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_78_446
timestamp 1
transform 1 0 41584 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_477
timestamp 1
transform 1 0 44436 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_483
timestamp 1
transform 1 0 44988 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_526
timestamp 1
transform 1 0 48944 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_78_533
timestamp 1
transform 1 0 49588 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_541
timestamp 1
transform 1 0 50324 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_584
timestamp 1
transform 1 0 54280 0 1 42976
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1636968456
transform 1 0 54740 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1636968456
transform 1 0 55844 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_613
timestamp 1636968456
transform 1 0 56948 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_625
timestamp 1636968456
transform 1 0 58052 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_637
timestamp 1
transform 1 0 59156 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_643
timestamp 1
transform 1 0 59708 0 1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_645
timestamp 1636968456
transform 1 0 59892 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_657
timestamp 1636968456
transform 1 0 60996 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_669
timestamp 1636968456
transform 1 0 62100 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_681
timestamp 1636968456
transform 1 0 63204 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_693
timestamp 1
transform 1 0 64308 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_699
timestamp 1
transform 1 0 64860 0 1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_701
timestamp 1636968456
transform 1 0 65044 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1636968456
transform 1 0 828 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1636968456
transform 1 0 1932 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1636968456
transform 1 0 3036 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1636968456
transform 1 0 4140 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1
transform 1 0 5244 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1
transform 1 0 5612 0 -1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1636968456
transform 1 0 5796 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1636968456
transform 1 0 6900 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1636968456
transform 1 0 8004 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1636968456
transform 1 0 9108 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1
transform 1 0 10212 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1
transform 1 0 10764 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_113
timestamp 1
transform 1 0 10948 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_169
timestamp 1
transform 1 0 16100 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_191
timestamp 1
transform 1 0 18124 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_225
timestamp 1
transform 1 0 21252 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_275
timestamp 1
transform 1 0 25852 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_289
timestamp 1
transform 1 0 27140 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_334
timestamp 1
transform 1 0 31280 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_337
timestamp 1
transform 1 0 31556 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_382
timestamp 1
transform 1 0 35696 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_421
timestamp 1
transform 1 0 39284 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1
transform 1 0 41676 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_479
timestamp 1
transform 1 0 44620 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_483
timestamp 1
transform 1 0 44988 0 -1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_522
timestamp 1636968456
transform 1 0 48576 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_534
timestamp 1636968456
transform 1 0 49680 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_546
timestamp 1636968456
transform 1 0 50784 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_558
timestamp 1
transform 1 0 51888 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_571
timestamp 1
transform 1 0 53084 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_575
timestamp 1
transform 1 0 53452 0 -1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_582
timestamp 1636968456
transform 1 0 54096 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_594
timestamp 1636968456
transform 1 0 55200 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_606
timestamp 1
transform 1 0 56304 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_614
timestamp 1
transform 1 0 57040 0 -1 44064
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_617
timestamp 1636968456
transform 1 0 57316 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_629
timestamp 1636968456
transform 1 0 58420 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_641
timestamp 1636968456
transform 1 0 59524 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_653
timestamp 1636968456
transform 1 0 60628 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_665
timestamp 1
transform 1 0 61732 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_671
timestamp 1
transform 1 0 62284 0 -1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_673
timestamp 1636968456
transform 1 0 62468 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_685
timestamp 1636968456
transform 1 0 63572 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_697
timestamp 1636968456
transform 1 0 64676 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_709
timestamp 1
transform 1 0 65780 0 -1 44064
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1636968456
transform 1 0 828 0 1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1636968456
transform 1 0 1932 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1
transform 1 0 3036 0 1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1636968456
transform 1 0 3220 0 1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1636968456
transform 1 0 4324 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_53
timestamp 1
transform 1 0 5428 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_57
timestamp 1
transform 1 0 5796 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_80_64
timestamp 1
transform 1 0 6440 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_80_70
timestamp 1
transform 1 0 6992 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_80_76
timestamp 1
transform 1 0 7544 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_80_82
timestamp 1
transform 1 0 8096 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_80_88
timestamp 1
transform 1 0 8648 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_80_94
timestamp 1
transform 1 0 9200 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_80_100
timestamp 1
transform 1 0 9752 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_80_141
timestamp 1
transform 1 0 13524 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_80_169
timestamp 1
transform 1 0 16100 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_80_215
timestamp 1
transform 1 0 20332 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_80_225
timestamp 1
transform 1 0 21252 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_80_237
timestamp 1
transform 1 0 22356 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_253
timestamp 1
transform 1 0 23828 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_267
timestamp 1
transform 1 0 25116 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_287
timestamp 1
transform 1 0 26956 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_349
timestamp 1
transform 1 0 32660 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_373
timestamp 1
transform 1 0 34868 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_388
timestamp 1
transform 1 0 36248 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_80_410
timestamp 1
transform 1 0 38272 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1
transform 1 0 39100 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_427
timestamp 1
transform 1 0 39836 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_474
timestamp 1
transform 1 0 44160 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_483
timestamp 1
transform 1 0 44988 0 1 44064
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_511
timestamp 1636968456
transform 1 0 47564 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_523
timestamp 1
transform 1 0 48668 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1
transform 1 0 49404 0 1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1636968456
transform 1 0 49588 0 1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1636968456
transform 1 0 50692 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_557
timestamp 1
transform 1 0 51796 0 1 44064
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_561
timestamp 1636968456
transform 1 0 52164 0 1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_573
timestamp 1636968456
transform 1 0 53268 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_585
timestamp 1
transform 1 0 54372 0 1 44064
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1636968456
transform 1 0 54740 0 1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1636968456
transform 1 0 55844 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_613
timestamp 1
transform 1 0 56948 0 1 44064
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_617
timestamp 1636968456
transform 1 0 57316 0 1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_629
timestamp 1636968456
transform 1 0 58420 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_641
timestamp 1
transform 1 0 59524 0 1 44064
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_645
timestamp 1636968456
transform 1 0 59892 0 1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_657
timestamp 1636968456
transform 1 0 60996 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_669
timestamp 1
transform 1 0 62100 0 1 44064
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_673
timestamp 1636968456
transform 1 0 62468 0 1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_685
timestamp 1636968456
transform 1 0 63572 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_697
timestamp 1
transform 1 0 64676 0 1 44064
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_701
timestamp 1636968456
transform 1 0 65044 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform 1 0 28980 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform 1 0 29716 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform -1 0 27784 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform 1 0 21252 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform 1 0 25576 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1
transform 1 0 23000 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1
transform -1 0 66148 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1
transform -1 0 23368 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1
transform 1 0 19412 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1
transform 1 0 18584 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1
transform -1 0 51612 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1
transform 1 0 47012 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1
transform -1 0 35696 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1
transform 1 0 63388 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1
transform -1 0 66148 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1
transform -1 0 66148 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1
transform -1 0 29072 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1
transform 1 0 14444 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1
transform -1 0 66148 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1
transform 1 0 17112 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1
transform 1 0 14444 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1
transform -1 0 17112 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1
transform -1 0 66148 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1
transform -1 0 66148 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1
transform -1 0 66148 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1
transform -1 0 66148 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1
transform -1 0 14076 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1
transform -1 0 27140 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1
transform -1 0 32016 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1
transform -1 0 34040 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1
transform -1 0 53176 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1
transform -1 0 51336 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1
transform -1 0 12696 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1
transform -1 0 29716 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1
transform -1 0 31464 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1
transform -1 0 16192 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1
transform -1 0 46368 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1
transform -1 0 8280 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1
transform -1 0 24564 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1
transform 1 0 37536 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1
transform 1 0 12696 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1
transform -1 0 53912 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1
transform -1 0 9752 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1
transform -1 0 57132 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1
transform -1 0 41768 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1
transform -1 0 53728 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1
transform -1 0 44068 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1
transform -1 0 40664 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1
transform -1 0 27876 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1
transform -1 0 66148 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1
transform 1 0 7544 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1
transform -1 0 9660 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1
transform -1 0 66148 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1
transform -1 0 54464 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1
transform 1 0 31556 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1
transform -1 0 35604 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1
transform -1 0 47380 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1
transform -1 0 66148 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1
transform -1 0 56672 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1
transform -1 0 65872 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1
transform -1 0 49404 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1
transform -1 0 52900 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1
transform -1 0 49496 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1
transform -1 0 61088 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1
transform -1 0 34868 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1
transform 1 0 38456 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1
transform -1 0 46000 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1
transform -1 0 66148 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1
transform 1 0 48392 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1
transform -1 0 64584 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1
transform -1 0 12604 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1
transform -1 0 21896 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1
transform -1 0 16008 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1
transform 1 0 23276 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1
transform 1 0 20424 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1
transform -1 0 38272 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1
transform 1 0 17848 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1
transform 1 0 65412 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1
transform -1 0 34868 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1
transform -1 0 19320 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1
transform -1 0 23736 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1
transform -1 0 45264 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1
transform -1 0 31188 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1
transform 1 0 15272 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1
transform -1 0 60628 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1
transform -1 0 41952 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1
transform -1 0 29808 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1
transform 1 0 47840 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1
transform -1 0 29808 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1
transform -1 0 66148 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1
transform 1 0 22080 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1
transform -1 0 44160 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1
transform -1 0 66148 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1
transform -1 0 66148 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1
transform -1 0 23276 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1
transform 1 0 13708 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1
transform 1 0 37812 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1
transform 1 0 14444 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1
transform -1 0 39284 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1
transform -1 0 46920 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1
transform -1 0 43424 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1
transform -1 0 34868 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1
transform 1 0 35052 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1
transform 1 0 32200 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1
transform -1 0 39008 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1
transform -1 0 32292 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1
transform -1 0 29992 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1
transform -1 0 30544 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1
transform -1 0 27140 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1
transform -1 0 33120 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1
transform 1 0 34132 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1
transform -1 0 27140 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1
transform 1 0 31188 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1
transform 1 0 27784 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1
transform -1 0 24288 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1
transform 1 0 26404 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_2_Left_66
timestamp 1
transform 1 0 63572 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_2_Right_147
timestamp 1
transform -1 0 66424 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_2_Left_0
timestamp 1
transform 1 0 63572 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_2_Right_67
timestamp 1
transform -1 0 66424 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_2_Left_1
timestamp 1
transform 1 0 63572 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_2_Right_68
timestamp 1
transform -1 0 66424 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_2_Left_2
timestamp 1
transform 1 0 63572 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_2_Right_69
timestamp 1
transform -1 0 66424 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_2_Left_3
timestamp 1
transform 1 0 63572 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_2_Right_70
timestamp 1
transform -1 0 66424 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_2_Left_4
timestamp 1
transform 1 0 63572 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_2_Right_71
timestamp 1
transform -1 0 66424 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_2_Left_5
timestamp 1
transform 1 0 63572 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_2_Right_72
timestamp 1
transform -1 0 66424 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_2_Left_6
timestamp 1
transform 1 0 63572 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_2_Right_73
timestamp 1
transform -1 0 66424 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_2_Left_7
timestamp 1
transform 1 0 63572 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_2_Right_74
timestamp 1
transform -1 0 66424 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_2_Left_8
timestamp 1
transform 1 0 63572 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_2_Right_75
timestamp 1
transform -1 0 66424 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Left_9
timestamp 1
transform 1 0 63572 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Right_76
timestamp 1
transform -1 0 66424 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Left_10
timestamp 1
transform 1 0 63572 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Right_77
timestamp 1
transform -1 0 66424 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Left_11
timestamp 1
transform 1 0 63572 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Right_78
timestamp 1
transform -1 0 66424 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Left_12
timestamp 1
transform 1 0 63572 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Right_79
timestamp 1
transform -1 0 66424 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Left_13
timestamp 1
transform 1 0 63572 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Right_80
timestamp 1
transform -1 0 66424 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Left_14
timestamp 1
transform 1 0 63572 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Right_81
timestamp 1
transform -1 0 66424 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Left_15
timestamp 1
transform 1 0 63572 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Right_82
timestamp 1
transform -1 0 66424 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Left_16
timestamp 1
transform 1 0 63572 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Right_83
timestamp 1
transform -1 0 66424 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Left_17
timestamp 1
transform 1 0 63572 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Right_84
timestamp 1
transform -1 0 66424 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Left_18
timestamp 1
transform 1 0 63572 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Right_85
timestamp 1
transform -1 0 66424 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Left_19
timestamp 1
transform 1 0 63572 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Right_86
timestamp 1
transform -1 0 66424 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Left_20
timestamp 1
transform 1 0 63572 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Right_87
timestamp 1
transform -1 0 66424 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Left_21
timestamp 1
transform 1 0 63572 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Right_88
timestamp 1
transform -1 0 66424 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Left_22
timestamp 1
transform 1 0 63572 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Right_89
timestamp 1
transform -1 0 66424 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Left_23
timestamp 1
transform 1 0 63572 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Right_90
timestamp 1
transform -1 0 66424 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Left_24
timestamp 1
transform 1 0 63572 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Right_91
timestamp 1
transform -1 0 66424 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Left_25
timestamp 1
transform 1 0 63572 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Right_92
timestamp 1
transform -1 0 66424 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Left_26
timestamp 1
transform 1 0 63572 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Right_93
timestamp 1
transform -1 0 66424 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Left_27
timestamp 1
transform 1 0 63572 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Right_94
timestamp 1
transform -1 0 66424 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Left_28
timestamp 1
transform 1 0 63572 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Right_95
timestamp 1
transform -1 0 66424 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Left_29
timestamp 1
transform 1 0 63572 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Right_96
timestamp 1
transform -1 0 66424 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Left_30
timestamp 1
transform 1 0 63572 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Right_97
timestamp 1
transform -1 0 66424 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Left_31
timestamp 1
transform 1 0 63572 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Right_98
timestamp 1
transform -1 0 66424 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Left_32
timestamp 1
transform 1 0 63572 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Right_99
timestamp 1
transform -1 0 66424 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Left_33
timestamp 1
transform 1 0 63572 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Right_100
timestamp 1
transform -1 0 66424 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Left_34
timestamp 1
transform 1 0 63572 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Right_101
timestamp 1
transform -1 0 66424 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Left_35
timestamp 1
transform 1 0 63572 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Right_102
timestamp 1
transform -1 0 66424 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Left_36
timestamp 1
transform 1 0 63572 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Right_103
timestamp 1
transform -1 0 66424 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Left_37
timestamp 1
transform 1 0 63572 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Right_104
timestamp 1
transform -1 0 66424 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Left_38
timestamp 1
transform 1 0 63572 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Right_105
timestamp 1
transform -1 0 66424 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Left_39
timestamp 1
transform 1 0 63572 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Right_106
timestamp 1
transform -1 0 66424 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Left_40
timestamp 1
transform 1 0 63572 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Right_107
timestamp 1
transform -1 0 66424 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Left_41
timestamp 1
transform 1 0 63572 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Right_108
timestamp 1
transform -1 0 66424 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Left_42
timestamp 1
transform 1 0 63572 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Right_109
timestamp 1
transform -1 0 66424 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Left_43
timestamp 1
transform 1 0 63572 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Right_110
timestamp 1
transform -1 0 66424 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Left_44
timestamp 1
transform 1 0 63572 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Right_111
timestamp 1
transform -1 0 66424 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Left_45
timestamp 1
transform 1 0 63572 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Right_112
timestamp 1
transform -1 0 66424 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Left_46
timestamp 1
transform 1 0 63572 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Right_113
timestamp 1
transform -1 0 66424 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Left_47
timestamp 1
transform 1 0 63572 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Right_114
timestamp 1
transform -1 0 66424 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Left_48
timestamp 1
transform 1 0 63572 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Right_115
timestamp 1
transform -1 0 66424 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Left_49
timestamp 1
transform 1 0 63572 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Right_116
timestamp 1
transform -1 0 66424 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Left_50
timestamp 1
transform 1 0 63572 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Right_117
timestamp 1
transform -1 0 66424 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Left_51
timestamp 1
transform 1 0 63572 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Right_118
timestamp 1
transform -1 0 66424 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Left_52
timestamp 1
transform 1 0 63572 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Right_119
timestamp 1
transform -1 0 66424 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Left_53
timestamp 1
transform 1 0 63572 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Right_120
timestamp 1
transform -1 0 66424 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Left_54
timestamp 1
transform 1 0 63572 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Right_121
timestamp 1
transform -1 0 66424 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Left_55
timestamp 1
transform 1 0 63572 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Right_122
timestamp 1
transform -1 0 66424 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Left_56
timestamp 1
transform 1 0 63572 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Right_123
timestamp 1
transform -1 0 66424 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Left_57
timestamp 1
transform 1 0 63572 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Right_124
timestamp 1
transform -1 0 66424 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Left_58
timestamp 1
transform 1 0 63572 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Right_125
timestamp 1
transform -1 0 66424 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Left_59
timestamp 1
transform 1 0 63572 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Right_126
timestamp 1
transform -1 0 66424 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Left_60
timestamp 1
transform 1 0 63572 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Right_127
timestamp 1
transform -1 0 66424 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Left_61
timestamp 1
transform 1 0 63572 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Right_128
timestamp 1
transform -1 0 66424 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Left_62
timestamp 1
transform 1 0 63572 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Right_129
timestamp 1
transform -1 0 66424 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Left_63
timestamp 1
transform 1 0 63572 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Right_130
timestamp 1
transform -1 0 66424 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Left_64
timestamp 1
transform 1 0 63572 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Right_131
timestamp 1
transform -1 0 66424 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Left_65
timestamp 1
transform 1 0 63572 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Right_132
timestamp 1
transform -1 0 66424 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_148
timestamp 1
transform 1 0 552 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_133
timestamp 1
transform -1 0 66424 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_149
timestamp 1
transform 1 0 552 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_134
timestamp 1
transform -1 0 66424 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Left_150
timestamp 1
transform 1 0 552 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Right_135
timestamp 1
transform -1 0 66424 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Left_151
timestamp 1
transform 1 0 552 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Right_136
timestamp 1
transform -1 0 66424 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Left_152
timestamp 1
transform 1 0 552 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Right_137
timestamp 1
transform -1 0 66424 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Left_153
timestamp 1
transform 1 0 552 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Right_138
timestamp 1
transform -1 0 66424 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Left_154
timestamp 1
transform 1 0 552 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Right_139
timestamp 1
transform -1 0 66424 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Left_155
timestamp 1
transform 1 0 552 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Right_140
timestamp 1
transform -1 0 66424 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Left_156
timestamp 1
transform 1 0 552 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Right_141
timestamp 1
transform -1 0 66424 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Left_157
timestamp 1
transform 1 0 552 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Right_142
timestamp 1
transform -1 0 66424 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Left_158
timestamp 1
transform 1 0 552 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Right_143
timestamp 1
transform -1 0 66424 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Left_159
timestamp 1
transform 1 0 552 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Right_144
timestamp 1
transform -1 0 66424 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Left_160
timestamp 1
transform 1 0 552 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Right_145
timestamp 1
transform -1 0 66424 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Left_161
timestamp 1
transform 1 0 552 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Right_146
timestamp 1
transform -1 0 66424 0 1 44064
box -38 -48 314 592
use sky130_sram_128B_1rw_32x32  SRAM
timestamp 0
transform -1 0 62536 0 -1 35514
box 0 0 1 1
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_162
timestamp 1
transform 1 0 3128 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_163
timestamp 1
transform 1 0 5704 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_164
timestamp 1
transform 1 0 8280 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_165
timestamp 1
transform 1 0 10856 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_166
timestamp 1
transform 1 0 13432 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_167
timestamp 1
transform 1 0 16008 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_168
timestamp 1
transform 1 0 18584 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_169
timestamp 1
transform 1 0 21160 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_170
timestamp 1
transform 1 0 23736 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_171
timestamp 1
transform 1 0 26312 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_172
timestamp 1
transform 1 0 28888 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_173
timestamp 1
transform 1 0 31464 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_174
timestamp 1
transform 1 0 34040 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_175
timestamp 1
transform 1 0 36616 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_176
timestamp 1
transform 1 0 39192 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_177
timestamp 1
transform 1 0 41768 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_178
timestamp 1
transform 1 0 44344 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_179
timestamp 1
transform 1 0 46920 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_180
timestamp 1
transform 1 0 49496 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_181
timestamp 1
transform 1 0 52072 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_182
timestamp 1
transform 1 0 54648 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_183
timestamp 1
transform 1 0 57224 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_184
timestamp 1
transform 1 0 59800 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_185
timestamp 1
transform 1 0 62376 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_186
timestamp 1
transform 1 0 64952 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_187
timestamp 1
transform 1 0 3128 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_188
timestamp 1
transform 1 0 8280 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_189
timestamp 1
transform 1 0 13432 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_190
timestamp 1
transform 1 0 18584 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_191
timestamp 1
transform 1 0 23736 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_192
timestamp 1
transform 1 0 28888 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_193
timestamp 1
transform 1 0 34040 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_194
timestamp 1
transform 1 0 39192 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_195
timestamp 1
transform 1 0 44344 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_196
timestamp 1
transform 1 0 49496 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_197
timestamp 1
transform 1 0 54648 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_198
timestamp 1
transform 1 0 59800 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_199
timestamp 1
transform 1 0 64952 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_200
timestamp 1
transform 1 0 5704 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_201
timestamp 1
transform 1 0 10856 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_202
timestamp 1
transform 1 0 16008 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_203
timestamp 1
transform 1 0 21160 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_204
timestamp 1
transform 1 0 26312 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_205
timestamp 1
transform 1 0 31464 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_206
timestamp 1
transform 1 0 36616 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_207
timestamp 1
transform 1 0 41768 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_208
timestamp 1
transform 1 0 46920 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_209
timestamp 1
transform 1 0 52072 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_210
timestamp 1
transform 1 0 57224 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_211
timestamp 1
transform 1 0 62376 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_212
timestamp 1
transform 1 0 3128 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_213
timestamp 1
transform 1 0 8280 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_214
timestamp 1
transform 1 0 13432 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_215
timestamp 1
transform 1 0 18584 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_216
timestamp 1
transform 1 0 23736 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_217
timestamp 1
transform 1 0 28888 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_218
timestamp 1
transform 1 0 34040 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_219
timestamp 1
transform 1 0 39192 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_220
timestamp 1
transform 1 0 44344 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_221
timestamp 1
transform 1 0 49496 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_222
timestamp 1
transform 1 0 54648 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_223
timestamp 1
transform 1 0 59800 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_224
timestamp 1
transform 1 0 64952 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_225
timestamp 1
transform 1 0 5704 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_226
timestamp 1
transform 1 0 10856 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_227
timestamp 1
transform 1 0 16008 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_228
timestamp 1
transform 1 0 21160 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_229
timestamp 1
transform 1 0 26312 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_230
timestamp 1
transform 1 0 31464 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_231
timestamp 1
transform 1 0 36616 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_232
timestamp 1
transform 1 0 41768 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_233
timestamp 1
transform 1 0 46920 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_234
timestamp 1
transform 1 0 52072 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_235
timestamp 1
transform 1 0 57224 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_236
timestamp 1
transform 1 0 62376 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_237
timestamp 1
transform 1 0 3128 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_238
timestamp 1
transform 1 0 8280 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_239
timestamp 1
transform 1 0 13432 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_240
timestamp 1
transform 1 0 18584 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_241
timestamp 1
transform 1 0 23736 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_242
timestamp 1
transform 1 0 28888 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_243
timestamp 1
transform 1 0 34040 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_244
timestamp 1
transform 1 0 39192 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_245
timestamp 1
transform 1 0 44344 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_246
timestamp 1
transform 1 0 49496 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_247
timestamp 1
transform 1 0 54648 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_248
timestamp 1
transform 1 0 59800 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_249
timestamp 1
transform 1 0 64952 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_250
timestamp 1
transform 1 0 5704 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_251
timestamp 1
transform 1 0 10856 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_252
timestamp 1
transform 1 0 16008 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_253
timestamp 1
transform 1 0 21160 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_254
timestamp 1
transform 1 0 26312 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_255
timestamp 1
transform 1 0 31464 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_256
timestamp 1
transform 1 0 36616 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_257
timestamp 1
transform 1 0 41768 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_258
timestamp 1
transform 1 0 46920 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_259
timestamp 1
transform 1 0 52072 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_260
timestamp 1
transform 1 0 57224 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_261
timestamp 1
transform 1 0 62376 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_262
timestamp 1
transform 1 0 3128 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_263
timestamp 1
transform 1 0 8280 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_264
timestamp 1
transform 1 0 13432 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_265
timestamp 1
transform 1 0 18584 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_266
timestamp 1
transform 1 0 23736 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_267
timestamp 1
transform 1 0 28888 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_268
timestamp 1
transform 1 0 34040 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_269
timestamp 1
transform 1 0 39192 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_270
timestamp 1
transform 1 0 44344 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_271
timestamp 1
transform 1 0 49496 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_272
timestamp 1
transform 1 0 54648 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_273
timestamp 1
transform 1 0 59800 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_274
timestamp 1
transform 1 0 64952 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_275
timestamp 1
transform 1 0 5704 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_276
timestamp 1
transform 1 0 10856 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_277
timestamp 1
transform 1 0 16008 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_278
timestamp 1
transform 1 0 21160 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_279
timestamp 1
transform 1 0 26312 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_280
timestamp 1
transform 1 0 31464 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_281
timestamp 1
transform 1 0 36616 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_282
timestamp 1
transform 1 0 41768 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_283
timestamp 1
transform 1 0 46920 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_284
timestamp 1
transform 1 0 52072 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_285
timestamp 1
transform 1 0 57224 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_286
timestamp 1
transform 1 0 62376 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_287
timestamp 1
transform 1 0 3128 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_288
timestamp 1
transform 1 0 8280 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_289
timestamp 1
transform 1 0 13432 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_290
timestamp 1
transform 1 0 18584 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_291
timestamp 1
transform 1 0 23736 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_292
timestamp 1
transform 1 0 28888 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_293
timestamp 1
transform 1 0 34040 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_294
timestamp 1
transform 1 0 39192 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_295
timestamp 1
transform 1 0 44344 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_296
timestamp 1
transform 1 0 49496 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_297
timestamp 1
transform 1 0 54648 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_298
timestamp 1
transform 1 0 59800 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_299
timestamp 1
transform 1 0 64952 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_300
timestamp 1
transform 1 0 5704 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_301
timestamp 1
transform 1 0 10856 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_302
timestamp 1
transform 1 0 16008 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_303
timestamp 1
transform 1 0 21160 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_304
timestamp 1
transform 1 0 26312 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_305
timestamp 1
transform 1 0 31464 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_306
timestamp 1
transform 1 0 36616 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_307
timestamp 1
transform 1 0 41768 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_308
timestamp 1
transform 1 0 46920 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_309
timestamp 1
transform 1 0 52072 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_310
timestamp 1
transform 1 0 57224 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_311
timestamp 1
transform 1 0 62376 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_312
timestamp 1
transform 1 0 3128 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_313
timestamp 1
transform 1 0 8280 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_314
timestamp 1
transform 1 0 13432 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_315
timestamp 1
transform 1 0 18584 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_316
timestamp 1
transform 1 0 23736 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_317
timestamp 1
transform 1 0 28888 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_318
timestamp 1
transform 1 0 34040 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_319
timestamp 1
transform 1 0 39192 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_320
timestamp 1
transform 1 0 44344 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_321
timestamp 1
transform 1 0 49496 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_322
timestamp 1
transform 1 0 54648 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_323
timestamp 1
transform 1 0 59800 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_324
timestamp 1
transform 1 0 64952 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_325
timestamp 1
transform 1 0 5704 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_326
timestamp 1
transform 1 0 10856 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_327
timestamp 1
transform 1 0 16008 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_328
timestamp 1
transform 1 0 21160 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_329
timestamp 1
transform 1 0 26312 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_330
timestamp 1
transform 1 0 31464 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_331
timestamp 1
transform 1 0 36616 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_332
timestamp 1
transform 1 0 41768 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_333
timestamp 1
transform 1 0 46920 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_334
timestamp 1
transform 1 0 52072 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_335
timestamp 1
transform 1 0 57224 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_336
timestamp 1
transform 1 0 62376 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_337
timestamp 1
transform 1 0 3128 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_338
timestamp 1
transform 1 0 5704 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_339
timestamp 1
transform 1 0 8280 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_340
timestamp 1
transform 1 0 10856 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_341
timestamp 1
transform 1 0 13432 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_342
timestamp 1
transform 1 0 16008 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_343
timestamp 1
transform 1 0 18584 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_344
timestamp 1
transform 1 0 21160 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_345
timestamp 1
transform 1 0 23736 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_346
timestamp 1
transform 1 0 26312 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_347
timestamp 1
transform 1 0 28888 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_348
timestamp 1
transform 1 0 31464 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_349
timestamp 1
transform 1 0 34040 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_350
timestamp 1
transform 1 0 36616 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_351
timestamp 1
transform 1 0 39192 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_352
timestamp 1
transform 1 0 41768 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_353
timestamp 1
transform 1 0 44344 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_354
timestamp 1
transform 1 0 46920 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_355
timestamp 1
transform 1 0 49496 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_356
timestamp 1
transform 1 0 52072 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_357
timestamp 1
transform 1 0 54648 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_358
timestamp 1
transform 1 0 57224 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_359
timestamp 1
transform 1 0 59800 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_360
timestamp 1
transform 1 0 62376 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_361
timestamp 1
transform 1 0 64952 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_57
timestamp 1
transform -1 0 10304 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_58
timestamp 1
transform -1 0 9752 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_59
timestamp 1
transform -1 0 9200 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_60
timestamp 1
transform -1 0 8648 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_61
timestamp 1
transform -1 0 8096 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_62
timestamp 1
transform -1 0 7544 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_63
timestamp 1
transform -1 0 6992 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_64
timestamp 1
transform -1 0 6440 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_65
timestamp 1
transform 1 0 12328 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_66
timestamp 1
transform 1 0 11776 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_67
timestamp 1
transform 1 0 11500 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_68
timestamp 1
transform 1 0 12604 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_69
timestamp 1
transform 1 0 11224 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_70
timestamp 1
transform 1 0 10948 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_71
timestamp 1
transform 1 0 10580 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_72
timestamp 1
transform 1 0 10304 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_73
timestamp 1
transform -1 0 20332 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_74
timestamp 1
transform -1 0 17756 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_75
timestamp 1
transform -1 0 17572 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_76
timestamp 1
transform -1 0 16468 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_77
timestamp 1
transform 1 0 12604 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_78
timestamp 1
transform 1 0 12052 0 1 44064
box -38 -48 314 592
<< labels >>
flabel metal4 s 2912 34210 3232 44656 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 50912 34142 51232 44656 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 65252 496 65572 37584 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1992 34208 2312 44656 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 49992 34142 50312 44656 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 64332 496 64652 37584 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 2 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 3 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 4 nsew signal input
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 5 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 6 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 7 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 8 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 9 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 10 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 11 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 12 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 13 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 14 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 15 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 16 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 17 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 18 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 19 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 20 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 21 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 22 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 23 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 24 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 25 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 26 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 27 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 28 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 29 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 30 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 31 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 32 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 33 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 34 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 35 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 36 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 37 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 38 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 39 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 40 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 41 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 42 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 43 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 44 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 66976 45152
<< end >>
