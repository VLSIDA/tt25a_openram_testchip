magic
tech sky130A
magscale 1 2
timestamp 1756846167
<< viali >>
rect 6193 44489 6227 44523
rect 6745 44489 6779 44523
rect 7297 44489 7331 44523
rect 7849 44489 7883 44523
rect 8401 44489 8435 44523
rect 8953 44489 8987 44523
rect 9505 44489 9539 44523
rect 10057 44489 10091 44523
rect 10609 44489 10643 44523
rect 12265 44489 12299 44523
rect 12541 44489 12575 44523
rect 12817 44489 12851 44523
rect 13553 44489 13587 44523
rect 13829 44489 13863 44523
rect 15485 44489 15519 44523
rect 15945 44489 15979 44523
rect 16221 44489 16255 44523
rect 16681 44489 16715 44523
rect 16957 44489 16991 44523
rect 17233 44489 17267 44523
rect 30849 44489 30883 44523
rect 40233 44489 40267 44523
rect 24961 44421 24995 44455
rect 30389 44421 30423 44455
rect 19349 44353 19383 44387
rect 20545 44353 20579 44387
rect 22477 44353 22511 44387
rect 25697 44353 25731 44387
rect 26801 44353 26835 44387
rect 27537 44353 27571 44387
rect 28825 44353 28859 44387
rect 33517 44353 33551 44387
rect 34989 44353 35023 44387
rect 37197 44353 37231 44387
rect 38025 44353 38059 44387
rect 42533 44353 42567 44387
rect 43269 44353 43303 44387
rect 46765 44353 46799 44387
rect 48145 44353 48179 44387
rect 10977 44285 11011 44319
rect 14657 44285 14691 44319
rect 17711 44285 17745 44319
rect 18521 44285 18555 44319
rect 20085 44285 20119 44319
rect 21097 44285 21131 44319
rect 22201 44285 22235 44319
rect 23489 44285 23523 44319
rect 24041 44285 24075 44319
rect 24409 44285 24443 44319
rect 26617 44285 26651 44319
rect 28273 44285 28307 44319
rect 30021 44285 30055 44319
rect 30757 44285 30791 44319
rect 31309 44285 31343 44319
rect 35817 44285 35851 44319
rect 36921 44285 36955 44319
rect 37841 44285 37875 44319
rect 38301 44285 38335 44319
rect 39681 44285 39715 44319
rect 40417 44285 40451 44319
rect 40969 44285 41003 44319
rect 44097 44285 44131 44319
rect 47593 44285 47627 44319
rect 11713 44217 11747 44251
rect 12081 44217 12115 44251
rect 14473 44217 14507 44251
rect 19073 44217 19107 44251
rect 19533 44217 19567 44251
rect 21281 44217 21315 44251
rect 21649 44217 21683 44251
rect 23857 44217 23891 44251
rect 25881 44217 25915 44251
rect 26065 44217 26099 44251
rect 29193 44217 29227 44251
rect 30205 44217 30239 44251
rect 34805 44217 34839 44251
rect 35265 44217 35299 44251
rect 37933 44217 37967 44251
rect 39313 44217 39347 44251
rect 39957 44217 39991 44251
rect 40693 44217 40727 44251
rect 41245 44217 41279 44251
rect 43085 44217 43119 44251
rect 43545 44217 43579 44251
rect 46489 44217 46523 44251
rect 47041 44217 47075 44251
rect 47869 44217 47903 44251
rect 11621 44149 11655 44183
rect 14381 44149 14415 44183
rect 15301 44149 15335 44183
rect 17417 44149 17451 44183
rect 17877 44149 17911 44183
rect 18705 44149 18739 44183
rect 19165 44149 19199 44183
rect 21833 44149 21867 44183
rect 22293 44149 22327 44183
rect 22937 44149 22971 44183
rect 25053 44149 25087 44183
rect 25421 44149 25455 44183
rect 25513 44149 25547 44183
rect 26433 44149 26467 44183
rect 27353 44149 27387 44183
rect 28089 44149 28123 44183
rect 29101 44149 29135 44183
rect 29377 44149 29411 44183
rect 31125 44149 31159 44183
rect 32965 44149 32999 44183
rect 33333 44149 33367 44183
rect 33425 44149 33459 44183
rect 34437 44149 34471 44183
rect 34897 44149 34931 44183
rect 37473 44149 37507 44183
rect 38945 44149 38979 44183
rect 41889 44149 41923 44183
rect 42257 44149 42291 44183
rect 42349 44149 42383 44183
rect 42717 44149 42751 44183
rect 43177 44149 43211 44183
rect 46121 44149 46155 44183
rect 46581 44149 46615 44183
rect 11989 43945 12023 43979
rect 14381 43945 14415 43979
rect 14841 43945 14875 43979
rect 19809 43945 19843 43979
rect 20269 43945 20303 43979
rect 36737 43945 36771 43979
rect 39773 43945 39807 43979
rect 43913 43945 43947 43979
rect 46857 43945 46891 43979
rect 47409 43945 47443 43979
rect 16497 43877 16531 43911
rect 17325 43877 17359 43911
rect 19073 43877 19107 43911
rect 21557 43877 21591 43911
rect 27353 43877 27387 43911
rect 29653 43877 29687 43911
rect 33977 43877 34011 43911
rect 38209 43877 38243 43911
rect 42349 43877 42383 43911
rect 45385 43877 45419 43911
rect 11161 43809 11195 43843
rect 12081 43809 12115 43843
rect 15301 43809 15335 43843
rect 15669 43809 15703 43843
rect 16589 43809 16623 43843
rect 19349 43809 19383 43843
rect 20821 43809 20855 43843
rect 23489 43809 23523 43843
rect 26249 43809 26283 43843
rect 27169 43809 27203 43843
rect 29377 43809 29411 43843
rect 31861 43809 31895 43843
rect 32781 43809 32815 43843
rect 33241 43809 33275 43843
rect 35909 43809 35943 43843
rect 38485 43809 38519 43843
rect 38945 43809 38979 43843
rect 39405 43809 39439 43843
rect 44465 43809 44499 43843
rect 48237 43809 48271 43843
rect 12265 43741 12299 43775
rect 12633 43741 12667 43775
rect 12909 43741 12943 43775
rect 14933 43741 14967 43775
rect 15025 43741 15059 43775
rect 16773 43741 16807 43775
rect 17049 43741 17083 43775
rect 19901 43741 19935 43775
rect 20085 43741 20119 43775
rect 21281 43741 21315 43775
rect 23029 43741 23063 43775
rect 23857 43741 23891 43775
rect 24501 43741 24535 43775
rect 25973 43741 26007 43775
rect 26985 43741 27019 43775
rect 27537 43741 27571 43775
rect 27813 43741 27847 43775
rect 29285 43741 29319 43775
rect 31401 43741 31435 43775
rect 32229 43741 32263 43775
rect 33057 43741 33091 43775
rect 33149 43741 33183 43775
rect 33701 43741 33735 43775
rect 35449 43741 35483 43775
rect 36001 43741 36035 43775
rect 36185 43741 36219 43775
rect 38669 43741 38703 43775
rect 38853 43741 38887 43775
rect 41245 43741 41279 43775
rect 41521 43741 41555 43775
rect 42073 43741 42107 43775
rect 43821 43741 43855 43775
rect 45109 43741 45143 43775
rect 47501 43741 47535 43775
rect 47593 43741 47627 43775
rect 48697 43741 48731 43775
rect 14473 43673 14507 43707
rect 16129 43673 16163 43707
rect 24409 43673 24443 43707
rect 35541 43673 35575 43707
rect 39589 43673 39623 43707
rect 11621 43605 11655 43639
rect 15853 43605 15887 43639
rect 17601 43605 17635 43639
rect 19441 43605 19475 43639
rect 23213 43605 23247 43639
rect 26433 43605 26467 43639
rect 31677 43605 31711 43639
rect 33609 43605 33643 43639
rect 39313 43605 39347 43639
rect 47041 43605 47075 43639
rect 47961 43605 47995 43639
rect 49249 43605 49283 43639
rect 15301 43401 15335 43435
rect 19809 43401 19843 43435
rect 21925 43401 21959 43435
rect 22109 43401 22143 43435
rect 23949 43401 23983 43435
rect 26065 43401 26099 43435
rect 28641 43401 28675 43435
rect 29009 43401 29043 43435
rect 29837 43401 29871 43435
rect 34161 43401 34195 43435
rect 36645 43401 36679 43435
rect 39313 43401 39347 43435
rect 40325 43401 40359 43435
rect 42809 43401 42843 43435
rect 18797 43333 18831 43367
rect 42717 43333 42751 43367
rect 11069 43265 11103 43299
rect 11345 43265 11379 43299
rect 11437 43265 11471 43299
rect 13553 43265 13587 43299
rect 19165 43265 19199 43299
rect 21649 43265 21683 43299
rect 22661 43265 22695 43299
rect 26617 43265 26651 43299
rect 27537 43265 27571 43299
rect 27629 43265 27663 43299
rect 29653 43265 29687 43299
rect 30389 43265 30423 43299
rect 33701 43265 33735 43299
rect 33977 43265 34011 43299
rect 34897 43265 34931 43299
rect 37197 43265 37231 43299
rect 37473 43265 37507 43299
rect 38945 43265 38979 43299
rect 40969 43265 41003 43299
rect 43269 43265 43303 43299
rect 43361 43265 43395 43299
rect 45017 43265 45051 43299
rect 45845 43265 45879 43299
rect 47317 43265 47351 43299
rect 47685 43265 47719 43299
rect 16037 43197 16071 43231
rect 16221 43197 16255 43231
rect 18981 43197 19015 43231
rect 19441 43197 19475 43231
rect 21741 43197 21775 43231
rect 22569 43197 22603 43231
rect 23581 43197 23615 43231
rect 24133 43197 24167 43231
rect 24225 43197 24259 43231
rect 26433 43197 26467 43231
rect 27445 43197 27479 43231
rect 28457 43197 28491 43231
rect 28825 43197 28859 43231
rect 29377 43197 29411 43231
rect 30739 43197 30773 43231
rect 31217 43197 31251 43231
rect 31585 43197 31619 43231
rect 34713 43197 34747 43231
rect 39865 43197 39899 43231
rect 40877 43197 40911 43231
rect 43729 43197 43763 43231
rect 47593 43197 47627 43231
rect 49433 43197 49467 43231
rect 51825 43197 51859 43231
rect 11713 43129 11747 43163
rect 13829 43129 13863 43163
rect 16497 43129 16531 43163
rect 19349 43129 19383 43163
rect 21373 43129 21407 43163
rect 22477 43129 22511 43163
rect 24501 43129 24535 43163
rect 27905 43129 27939 43163
rect 30205 43129 30239 43163
rect 35173 43129 35207 43163
rect 40417 43129 40451 43163
rect 41245 43129 41279 43163
rect 43177 43129 43211 43163
rect 44281 43129 44315 43163
rect 44833 43129 44867 43163
rect 49157 43129 49191 43163
rect 52377 43129 52411 43163
rect 9597 43061 9631 43095
rect 13185 43061 13219 43095
rect 15485 43061 15519 43095
rect 17969 43061 18003 43095
rect 19901 43061 19935 43095
rect 22937 43061 22971 43095
rect 25973 43061 26007 43095
rect 26525 43061 26559 43095
rect 27077 43061 27111 43095
rect 29469 43061 29503 43095
rect 30297 43061 30331 43095
rect 30849 43061 30883 43095
rect 32229 43061 32263 43095
rect 40693 43061 40727 43095
rect 44465 43061 44499 43095
rect 44925 43061 44959 43095
rect 51273 43061 51307 43095
rect 52101 43061 52135 43095
rect 12081 42857 12115 42891
rect 12449 42857 12483 42891
rect 12909 42857 12943 42891
rect 13369 42857 13403 42891
rect 14105 42857 14139 42891
rect 20269 42857 20303 42891
rect 20729 42857 20763 42891
rect 22017 42857 22051 42891
rect 22753 42857 22787 42891
rect 24869 42857 24903 42891
rect 25789 42857 25823 42891
rect 26249 42857 26283 42891
rect 38669 42857 38703 42891
rect 39037 42857 39071 42891
rect 39129 42857 39163 42891
rect 40325 42857 40359 42891
rect 41061 42857 41095 42891
rect 41429 42857 41463 42891
rect 44373 42857 44407 42891
rect 44741 42857 44775 42891
rect 46581 42857 46615 42891
rect 47041 42857 47075 42891
rect 47409 42857 47443 42891
rect 48605 42857 48639 42891
rect 49065 42857 49099 42891
rect 49433 42857 49467 42891
rect 21649 42789 21683 42823
rect 27261 42789 27295 42823
rect 27353 42789 27387 42823
rect 28089 42789 28123 42823
rect 29377 42789 29411 42823
rect 30573 42789 30607 42823
rect 32413 42789 32447 42823
rect 34345 42789 34379 42823
rect 35357 42789 35391 42823
rect 37381 42789 37415 42823
rect 38209 42789 38243 42823
rect 39497 42789 39531 42823
rect 12541 42721 12575 42755
rect 13277 42721 13311 42755
rect 14749 42721 14783 42755
rect 15209 42721 15243 42755
rect 16129 42721 16163 42755
rect 18429 42721 18463 42755
rect 20637 42721 20671 42755
rect 22661 42721 22695 42755
rect 25881 42721 25915 42755
rect 26433 42721 26467 42755
rect 28825 42721 28859 42755
rect 29285 42721 29319 42755
rect 30665 42721 30699 42755
rect 35449 42721 35483 42755
rect 36553 42721 36587 42755
rect 36829 42721 36863 42755
rect 37289 42721 37323 42755
rect 38301 42721 38335 42755
rect 40509 42721 40543 42755
rect 42165 42721 42199 42755
rect 44925 42721 44959 42755
rect 46489 42721 46523 42755
rect 49985 42721 50019 42755
rect 52193 42721 52227 42755
rect 12725 42653 12759 42687
rect 13553 42653 13587 42687
rect 14197 42653 14231 42687
rect 14381 42653 14415 42687
rect 15393 42653 15427 42687
rect 16405 42653 16439 42687
rect 18705 42653 18739 42687
rect 20177 42653 20211 42687
rect 20821 42653 20855 42687
rect 21465 42653 21499 42687
rect 21557 42653 21591 42687
rect 22845 42653 22879 42687
rect 23121 42653 23155 42687
rect 23397 42653 23431 42687
rect 25697 42653 25731 42687
rect 27537 42653 27571 42687
rect 28181 42653 28215 42687
rect 28365 42653 28399 42687
rect 29101 42653 29135 42687
rect 30757 42653 30791 42687
rect 32137 42653 32171 42687
rect 34437 42653 34471 42687
rect 34529 42653 34563 42687
rect 35173 42653 35207 42687
rect 37197 42653 37231 42687
rect 38485 42653 38519 42687
rect 39221 42653 39255 42687
rect 40049 42653 40083 42687
rect 40877 42653 40911 42687
rect 40969 42653 41003 42687
rect 42441 42653 42475 42687
rect 44189 42653 44223 42687
rect 44281 42653 44315 42687
rect 45569 42653 45603 42687
rect 46305 42653 46339 42687
rect 47501 42653 47535 42687
rect 47685 42653 47719 42687
rect 48697 42653 48731 42687
rect 48881 42653 48915 42687
rect 49525 42653 49559 42687
rect 49617 42653 49651 42687
rect 50261 42653 50295 42687
rect 54125 42653 54159 42687
rect 13737 42585 13771 42619
rect 15025 42585 15059 42619
rect 22293 42585 22327 42619
rect 26617 42585 26651 42619
rect 27721 42585 27755 42619
rect 29745 42585 29779 42619
rect 30205 42585 30239 42619
rect 33977 42585 34011 42619
rect 37749 42585 37783 42619
rect 52377 42585 52411 42619
rect 14657 42517 14691 42551
rect 15945 42517 15979 42551
rect 17877 42517 17911 42551
rect 22201 42517 22235 42551
rect 26893 42517 26927 42551
rect 28641 42517 28675 42551
rect 33885 42517 33919 42551
rect 34989 42517 35023 42551
rect 35817 42517 35851 42551
rect 35909 42517 35943 42551
rect 37841 42517 37875 42551
rect 43913 42517 43947 42551
rect 45661 42517 45695 42551
rect 48237 42517 48271 42551
rect 51733 42517 51767 42551
rect 53573 42517 53607 42551
rect 10149 42313 10183 42347
rect 16497 42313 16531 42347
rect 16773 42313 16807 42347
rect 20545 42313 20579 42347
rect 24685 42313 24719 42347
rect 28641 42313 28675 42347
rect 29009 42313 29043 42347
rect 34161 42313 34195 42347
rect 35081 42313 35115 42347
rect 35265 42313 35299 42347
rect 37013 42313 37047 42347
rect 38945 42313 38979 42347
rect 42073 42313 42107 42347
rect 10241 42245 10275 42279
rect 19625 42245 19659 42279
rect 23857 42245 23891 42279
rect 25697 42245 25731 42279
rect 30481 42245 30515 42279
rect 43453 42245 43487 42279
rect 8677 42177 8711 42211
rect 10885 42177 10919 42211
rect 11621 42177 11655 42211
rect 14749 42177 14783 42211
rect 17417 42177 17451 42211
rect 18061 42177 18095 42211
rect 18245 42177 18279 42211
rect 19165 42177 19199 42211
rect 19257 42177 19291 42211
rect 23029 42177 23063 42211
rect 24409 42177 24443 42211
rect 25145 42177 25179 42211
rect 25329 42177 25363 42211
rect 26157 42177 26191 42211
rect 26249 42177 26283 42211
rect 26893 42177 26927 42211
rect 27169 42177 27203 42211
rect 33425 42177 33459 42211
rect 34621 42177 34655 42211
rect 34713 42177 34747 42211
rect 35725 42177 35759 42211
rect 35817 42177 35851 42211
rect 37473 42177 37507 42211
rect 40785 42177 40819 42211
rect 42625 42177 42659 42211
rect 44005 42177 44039 42211
rect 44925 42177 44959 42211
rect 45017 42177 45051 42211
rect 47317 42177 47351 42211
rect 47409 42177 47443 42211
rect 47685 42177 47719 42211
rect 49433 42177 49467 42211
rect 52653 42177 52687 42211
rect 53389 42177 53423 42211
rect 54217 42177 54251 42211
rect 8401 42109 8435 42143
rect 17141 42109 17175 42143
rect 19073 42109 19107 42143
rect 23305 42109 23339 42143
rect 24225 42109 24259 42143
rect 29561 42109 29595 42143
rect 32137 42109 32171 42143
rect 33793 42109 33827 42143
rect 33977 42109 34011 42143
rect 35633 42109 35667 42143
rect 36093 42109 36127 42143
rect 37197 42109 37231 42143
rect 39957 42109 39991 42143
rect 41705 42109 41739 42143
rect 42533 42109 42567 42143
rect 42993 42109 43027 42143
rect 43821 42109 43855 42143
rect 53113 42109 53147 42143
rect 53941 42109 53975 42143
rect 55045 42109 55079 42143
rect 10609 42041 10643 42075
rect 11069 42041 11103 42075
rect 15025 42041 15059 42075
rect 17233 42041 17267 42075
rect 21833 42041 21867 42075
rect 26065 42041 26099 42075
rect 30757 42041 30791 42075
rect 32689 42041 32723 42075
rect 40601 42041 40635 42075
rect 41061 42041 41095 42075
rect 41889 42041 41923 42075
rect 42441 42041 42475 42075
rect 43361 42041 43395 42075
rect 43913 42041 43947 42075
rect 45293 42041 45327 42075
rect 47041 42041 47075 42075
rect 50629 42041 50663 42075
rect 52377 42041 52411 42075
rect 10701 41973 10735 42007
rect 17601 41973 17635 42007
rect 17969 41973 18003 42007
rect 18705 41973 18739 42007
rect 22385 41973 22419 42007
rect 23213 41973 23247 42007
rect 23673 41973 23707 42007
rect 24317 41973 24351 42007
rect 25053 41973 25087 42007
rect 25605 41973 25639 42007
rect 30297 41973 30331 42007
rect 32781 41973 32815 42007
rect 33149 41973 33183 42007
rect 33241 41973 33275 42007
rect 34529 41973 34563 42007
rect 39313 41973 39347 42007
rect 40233 41973 40267 42007
rect 40693 41973 40727 42007
rect 44465 41973 44499 42007
rect 44833 41973 44867 42007
rect 45569 41973 45603 42007
rect 52745 41973 52779 42007
rect 53205 41973 53239 42007
rect 53573 41973 53607 42007
rect 54033 41973 54067 42007
rect 54861 41973 54895 42007
rect 10425 41769 10459 41803
rect 15209 41769 15243 41803
rect 15577 41769 15611 41803
rect 15669 41769 15703 41803
rect 16405 41769 16439 41803
rect 17233 41769 17267 41803
rect 17601 41769 17635 41803
rect 17693 41769 17727 41803
rect 28641 41769 28675 41803
rect 33701 41769 33735 41803
rect 37197 41769 37231 41803
rect 41337 41769 41371 41803
rect 42441 41769 42475 41803
rect 44741 41769 44775 41803
rect 47041 41769 47075 41803
rect 48973 41769 49007 41803
rect 49065 41769 49099 41803
rect 49433 41769 49467 41803
rect 50261 41769 50295 41803
rect 50629 41769 50663 41803
rect 16865 41701 16899 41735
rect 23121 41701 23155 41735
rect 25697 41701 25731 41735
rect 26709 41701 26743 41735
rect 29009 41701 29043 41735
rect 32229 41701 32263 41735
rect 37657 41701 37691 41735
rect 39405 41701 39439 41735
rect 43269 41701 43303 41735
rect 47501 41701 47535 41735
rect 48329 41701 48363 41735
rect 50721 41701 50755 41735
rect 52469 41701 52503 41735
rect 54125 41701 54159 41735
rect 10517 41633 10551 41667
rect 12725 41633 12759 41667
rect 13185 41633 13219 41667
rect 14289 41633 14323 41667
rect 16773 41633 16807 41667
rect 19533 41633 19567 41667
rect 20729 41633 20763 41667
rect 21281 41633 21315 41667
rect 23857 41633 23891 41667
rect 26433 41633 26467 41667
rect 30205 41633 30239 41667
rect 35081 41633 35115 41667
rect 39589 41633 39623 41667
rect 45109 41633 45143 41667
rect 47409 41633 47443 41667
rect 48237 41633 48271 41667
rect 51089 41633 51123 41667
rect 54493 41633 54527 41667
rect 57713 41633 57747 41667
rect 7941 41565 7975 41599
rect 8217 41565 8251 41599
rect 10609 41565 10643 41599
rect 12173 41565 12207 41599
rect 12817 41565 12851 41599
rect 12909 41565 12943 41599
rect 13829 41565 13863 41599
rect 15853 41565 15887 41599
rect 16957 41565 16991 41599
rect 17877 41565 17911 41599
rect 18613 41565 18647 41599
rect 18981 41565 19015 41599
rect 20269 41565 20303 41599
rect 20821 41565 20855 41599
rect 21005 41565 21039 41599
rect 21557 41565 21591 41599
rect 23029 41565 23063 41599
rect 23765 41565 23799 41599
rect 24133 41565 24167 41599
rect 25605 41565 25639 41599
rect 28181 41565 28215 41599
rect 29101 41565 29135 41599
rect 29193 41565 29227 41599
rect 31953 41565 31987 41599
rect 34253 41565 34287 41599
rect 36553 41565 36587 41599
rect 37013 41565 37047 41599
rect 37105 41565 37139 41599
rect 39865 41565 39899 41599
rect 42533 41565 42567 41599
rect 42717 41565 42751 41599
rect 42993 41565 43027 41599
rect 45385 41565 45419 41599
rect 46857 41565 46891 41599
rect 47593 41565 47627 41599
rect 48421 41565 48455 41599
rect 48789 41565 48823 41599
rect 50813 41565 50847 41599
rect 52193 41565 52227 41599
rect 56149 41565 56183 41599
rect 56425 41565 56459 41599
rect 57069 41565 57103 41599
rect 30389 41497 30423 41531
rect 35265 41497 35299 41531
rect 47869 41497 47903 41531
rect 53941 41497 53975 41531
rect 9689 41429 9723 41463
rect 10057 41429 10091 41463
rect 11621 41429 11655 41463
rect 12357 41429 12391 41463
rect 14197 41429 14231 41463
rect 18061 41429 18095 41463
rect 19625 41429 19659 41463
rect 20361 41429 20395 41463
rect 34897 41429 34931 41463
rect 35909 41429 35943 41463
rect 37565 41429 37599 41463
rect 42073 41429 42107 41463
rect 54677 41429 54711 41463
rect 56517 41429 56551 41463
rect 57621 41429 57655 41463
rect 16773 41225 16807 41259
rect 19901 41225 19935 41259
rect 21833 41225 21867 41259
rect 24133 41225 24167 41259
rect 25697 41225 25731 41259
rect 33885 41225 33919 41259
rect 37657 41225 37691 41259
rect 37841 41225 37875 41259
rect 39313 41225 39347 41259
rect 47869 41225 47903 41259
rect 48605 41225 48639 41259
rect 53021 41225 53055 41259
rect 21741 41157 21775 41191
rect 34161 41157 34195 41191
rect 9413 41089 9447 41123
rect 9689 41089 9723 41123
rect 11437 41089 11471 41123
rect 11621 41089 11655 41123
rect 13369 41089 13403 41123
rect 13737 41089 13771 41123
rect 17509 41089 17543 41123
rect 18429 41089 18463 41123
rect 19993 41089 20027 41123
rect 20269 41089 20303 41123
rect 22385 41089 22419 41123
rect 23121 41089 23155 41123
rect 24685 41089 24719 41123
rect 30481 41089 30515 41123
rect 31861 41089 31895 41123
rect 32137 41089 32171 41123
rect 32413 41089 32447 41123
rect 34713 41089 34747 41123
rect 35541 41089 35575 41123
rect 38301 41089 38335 41123
rect 38485 41089 38519 41123
rect 39773 41089 39807 41123
rect 39865 41089 39899 41123
rect 43177 41089 43211 41123
rect 46949 41089 46983 41123
rect 47317 41089 47351 41123
rect 47961 41089 47995 41123
rect 50261 41089 50295 41123
rect 53481 41089 53515 41123
rect 53665 41089 53699 41123
rect 53941 41089 53975 41123
rect 55873 41089 55907 41123
rect 56701 41089 56735 41123
rect 57529 41089 57563 41123
rect 9321 41021 9355 41055
rect 13921 41021 13955 41055
rect 15025 41021 15059 41055
rect 17233 41021 17267 41055
rect 19257 41021 19291 41055
rect 24593 41021 24627 41055
rect 26985 41021 27019 41055
rect 27077 41021 27111 41055
rect 28825 41021 28859 41055
rect 30665 41021 30699 41055
rect 31217 41021 31251 41055
rect 31677 41021 31711 41055
rect 34529 41021 34563 41055
rect 35357 41021 35391 41055
rect 38669 41021 38703 41055
rect 41981 41021 42015 41055
rect 51181 41021 51215 41055
rect 56517 41021 56551 41055
rect 57621 41021 57655 41055
rect 57805 41021 57839 41055
rect 11897 40953 11931 40987
rect 15301 40953 15335 40987
rect 35909 40953 35943 40987
rect 37565 40953 37599 40987
rect 41705 40953 41739 40987
rect 42993 40953 43027 40987
rect 43361 40953 43395 40987
rect 44465 40953 44499 40987
rect 46213 40953 46247 40987
rect 46765 40953 46799 40987
rect 47409 40953 47443 40987
rect 47501 40953 47535 40987
rect 50077 40953 50111 40987
rect 54217 40953 54251 40987
rect 54861 40953 54895 40987
rect 56609 40953 56643 40987
rect 57069 40953 57103 40987
rect 8677 40885 8711 40919
rect 13829 40885 13863 40919
rect 14289 40885 14323 40919
rect 16865 40885 16899 40919
rect 17325 40885 17359 40919
rect 17877 40885 17911 40919
rect 22201 40885 22235 40919
rect 22293 40885 22327 40919
rect 23673 40885 23707 40919
rect 24501 40885 24535 40919
rect 29837 40885 29871 40919
rect 31309 40885 31343 40919
rect 31769 40885 31803 40919
rect 34621 40885 34655 40919
rect 34989 40885 35023 40919
rect 35449 40885 35483 40919
rect 38209 40885 38243 40919
rect 39681 40885 39715 40919
rect 40233 40885 40267 40919
rect 42533 40885 42567 40919
rect 42901 40885 42935 40919
rect 46305 40885 46339 40919
rect 46673 40885 46707 40919
rect 49709 40885 49743 40919
rect 50169 40885 50203 40919
rect 52469 40885 52503 40919
rect 53389 40885 53423 40919
rect 54953 40885 54987 40919
rect 55321 40885 55355 40919
rect 55689 40885 55723 40919
rect 55781 40885 55815 40919
rect 56149 40885 56183 40919
rect 57161 40885 57195 40919
rect 10977 40681 11011 40715
rect 11345 40681 11379 40715
rect 15945 40681 15979 40715
rect 17325 40681 17359 40715
rect 17877 40681 17911 40715
rect 21281 40681 21315 40715
rect 22201 40681 22235 40715
rect 25513 40681 25547 40715
rect 26801 40681 26835 40715
rect 29101 40681 29135 40715
rect 31401 40681 31435 40715
rect 32505 40681 32539 40715
rect 32965 40681 32999 40715
rect 34161 40681 34195 40715
rect 34529 40681 34563 40715
rect 36553 40681 36587 40715
rect 51273 40681 51307 40715
rect 14105 40613 14139 40647
rect 15485 40613 15519 40647
rect 17233 40613 17267 40647
rect 23949 40613 23983 40647
rect 25881 40613 25915 40647
rect 27261 40613 27295 40647
rect 29929 40613 29963 40647
rect 35081 40613 35115 40647
rect 37657 40613 37691 40647
rect 41889 40613 41923 40647
rect 45937 40613 45971 40647
rect 47409 40613 47443 40647
rect 49433 40613 49467 40647
rect 51641 40613 51675 40647
rect 55229 40613 55263 40647
rect 10793 40545 10827 40579
rect 11437 40545 11471 40579
rect 14381 40545 14415 40579
rect 15577 40545 15611 40579
rect 18245 40545 18279 40579
rect 19073 40545 19107 40579
rect 21649 40545 21683 40579
rect 22845 40545 22879 40579
rect 25973 40545 26007 40579
rect 27813 40545 27847 40579
rect 28733 40545 28767 40579
rect 29193 40545 29227 40579
rect 31677 40545 31711 40579
rect 32597 40545 32631 40579
rect 33333 40545 33367 40579
rect 33425 40545 33459 40579
rect 34805 40545 34839 40579
rect 37381 40545 37415 40579
rect 39589 40545 39623 40579
rect 40693 40545 40727 40579
rect 41613 40545 41647 40579
rect 45477 40545 45511 40579
rect 47501 40545 47535 40579
rect 52469 40545 52503 40579
rect 54861 40545 54895 40579
rect 54953 40545 54987 40579
rect 8769 40477 8803 40511
rect 9045 40477 9079 40511
rect 11621 40477 11655 40511
rect 12357 40477 12391 40511
rect 14565 40477 14599 40511
rect 15393 40477 15427 40511
rect 17417 40477 17451 40511
rect 17785 40477 17819 40511
rect 18337 40477 18371 40511
rect 18429 40477 18463 40511
rect 19349 40477 19383 40511
rect 21741 40477 21775 40511
rect 21925 40477 21959 40511
rect 23581 40477 23615 40511
rect 23673 40477 23707 40511
rect 26065 40477 26099 40511
rect 26893 40477 26927 40511
rect 27077 40477 27111 40511
rect 29009 40477 29043 40511
rect 29653 40477 29687 40511
rect 32689 40477 32723 40511
rect 33609 40477 33643 40511
rect 33977 40477 34011 40511
rect 34069 40477 34103 40511
rect 39129 40477 39163 40511
rect 39681 40477 39715 40511
rect 39773 40477 39807 40511
rect 40785 40477 40819 40511
rect 40877 40477 40911 40511
rect 43729 40477 43763 40511
rect 45201 40477 45235 40511
rect 46029 40477 46063 40511
rect 46121 40477 46155 40511
rect 47593 40477 47627 40511
rect 48513 40477 48547 40511
rect 49157 40477 49191 40511
rect 51181 40477 51215 40511
rect 51733 40477 51767 40511
rect 51825 40477 51859 40511
rect 52837 40477 52871 40511
rect 54585 40477 54619 40511
rect 56977 40477 57011 40511
rect 40325 40409 40359 40443
rect 45569 40409 45603 40443
rect 47041 40409 47075 40443
rect 15117 40341 15151 40375
rect 16865 40341 16899 40375
rect 20821 40341 20855 40375
rect 22937 40341 22971 40375
rect 25421 40341 25455 40375
rect 26433 40341 26467 40375
rect 28089 40341 28123 40375
rect 29561 40341 29595 40375
rect 31953 40341 31987 40375
rect 32137 40341 32171 40375
rect 39221 40341 39255 40375
rect 43361 40341 43395 40375
rect 49065 40341 49099 40375
rect 52653 40341 52687 40375
rect 9505 40137 9539 40171
rect 16300 40137 16334 40171
rect 20563 40137 20597 40171
rect 20913 40137 20947 40171
rect 22109 40137 22143 40171
rect 24133 40137 24167 40171
rect 26721 40137 26755 40171
rect 28825 40137 28859 40171
rect 37644 40137 37678 40171
rect 46685 40137 46719 40171
rect 49617 40137 49651 40171
rect 56333 40137 56367 40171
rect 49433 40069 49467 40103
rect 9321 40001 9355 40035
rect 9965 40001 9999 40035
rect 10149 40001 10183 40035
rect 10885 40001 10919 40035
rect 11805 40001 11839 40035
rect 13093 40001 13127 40035
rect 13277 40001 13311 40035
rect 14197 40001 14231 40035
rect 14473 40001 14507 40035
rect 16037 40001 16071 40035
rect 17785 40001 17819 40035
rect 20821 40001 20855 40035
rect 21465 40001 21499 40035
rect 22569 40001 22603 40035
rect 22661 40001 22695 40035
rect 23489 40001 23523 40035
rect 24593 40001 24627 40035
rect 24777 40001 24811 40035
rect 27077 40001 27111 40035
rect 29653 40001 29687 40035
rect 29837 40001 29871 40035
rect 37105 40001 37139 40035
rect 37381 40001 37415 40035
rect 39129 40001 39163 40035
rect 39497 40001 39531 40035
rect 40141 40001 40175 40035
rect 44005 40001 44039 40035
rect 44189 40001 44223 40035
rect 46949 40001 46983 40035
rect 48881 40001 48915 40035
rect 51089 40001 51123 40035
rect 51365 40001 51399 40035
rect 55689 40001 55723 40035
rect 57805 40001 57839 40035
rect 58633 40001 58667 40035
rect 13001 39933 13035 39967
rect 21281 39933 21315 39967
rect 23305 39933 23339 39967
rect 24501 39933 24535 39967
rect 26985 39933 27019 39967
rect 39681 39933 39715 39967
rect 40693 39933 40727 39967
rect 40877 39933 40911 39967
rect 47133 39933 47167 39967
rect 48053 39933 48087 39967
rect 49065 39933 49099 39967
rect 52009 39933 52043 39967
rect 57713 39933 57747 39967
rect 9045 39865 9079 39899
rect 9137 39865 9171 39899
rect 11529 39865 11563 39899
rect 21373 39865 21407 39899
rect 22477 39865 22511 39899
rect 27353 39865 27387 39899
rect 29377 39865 29411 39899
rect 30113 39865 30147 39899
rect 36829 39865 36863 39899
rect 41153 39865 41187 39899
rect 43361 39865 43395 39899
rect 43913 39865 43947 39899
rect 55873 39865 55907 39899
rect 56977 39865 57011 39899
rect 57621 39865 57655 39899
rect 8677 39797 8711 39831
rect 9873 39797 9907 39831
rect 10333 39797 10367 39831
rect 10701 39797 10735 39831
rect 10793 39797 10827 39831
rect 11161 39797 11195 39831
rect 11621 39797 11655 39831
rect 12633 39797 12667 39831
rect 15945 39797 15979 39831
rect 17969 39797 18003 39831
rect 19073 39797 19107 39831
rect 22937 39797 22971 39831
rect 23397 39797 23431 39831
rect 25237 39797 25271 39831
rect 29009 39797 29043 39831
rect 29469 39797 29503 39831
rect 31585 39797 31619 39831
rect 32965 39797 32999 39831
rect 35357 39797 35391 39831
rect 39589 39797 39623 39831
rect 40049 39797 40083 39831
rect 42625 39797 42659 39831
rect 43545 39797 43579 39831
rect 45201 39797 45235 39831
rect 47777 39797 47811 39831
rect 48605 39797 48639 39831
rect 48973 39797 49007 39831
rect 55413 39797 55447 39831
rect 55965 39797 55999 39831
rect 57253 39797 57287 39831
rect 58081 39797 58115 39831
rect 58449 39797 58483 39831
rect 58541 39797 58575 39831
rect 15209 39593 15243 39627
rect 15577 39593 15611 39627
rect 15669 39593 15703 39627
rect 16313 39593 16347 39627
rect 16773 39593 16807 39627
rect 18245 39593 18279 39627
rect 18705 39593 18739 39627
rect 20085 39593 20119 39627
rect 26249 39593 26283 39627
rect 26433 39593 26467 39627
rect 26893 39593 26927 39627
rect 27721 39593 27755 39627
rect 28089 39593 28123 39627
rect 30389 39593 30423 39627
rect 33793 39593 33827 39627
rect 35633 39593 35667 39627
rect 36737 39593 36771 39627
rect 38393 39593 38427 39627
rect 40693 39593 40727 39627
rect 42165 39593 42199 39627
rect 42257 39593 42291 39627
rect 46673 39593 46707 39627
rect 47409 39593 47443 39627
rect 48421 39593 48455 39627
rect 50537 39593 50571 39627
rect 50997 39593 51031 39627
rect 51549 39593 51583 39627
rect 54861 39593 54895 39627
rect 55229 39593 55263 39627
rect 55321 39593 55355 39627
rect 59461 39593 59495 39627
rect 10149 39525 10183 39559
rect 14473 39525 14507 39559
rect 16221 39525 16255 39559
rect 16681 39525 16715 39559
rect 18797 39525 18831 39559
rect 21741 39525 21775 39559
rect 22753 39525 22787 39559
rect 24777 39525 24811 39559
rect 26801 39525 26835 39559
rect 28825 39525 28859 39559
rect 32229 39525 32263 39559
rect 36093 39525 36127 39559
rect 37105 39525 37139 39559
rect 39865 39525 39899 39559
rect 51457 39525 51491 39559
rect 53757 39525 53791 39559
rect 57621 39525 57655 39559
rect 10425 39457 10459 39491
rect 11345 39457 11379 39491
rect 11437 39457 11471 39491
rect 14381 39457 14415 39491
rect 17509 39457 17543 39491
rect 17601 39457 17635 39491
rect 18337 39457 18371 39491
rect 21649 39457 21683 39491
rect 22477 39457 22511 39491
rect 24501 39457 24535 39491
rect 27445 39457 27479 39491
rect 30757 39457 30791 39491
rect 31953 39457 31987 39491
rect 34345 39457 34379 39491
rect 36001 39457 36035 39491
rect 40141 39457 40175 39491
rect 40601 39457 40635 39491
rect 43085 39457 43119 39491
rect 44925 39457 44959 39491
rect 50629 39457 50663 39491
rect 52193 39457 52227 39491
rect 54401 39457 54435 39491
rect 55689 39457 55723 39491
rect 8401 39389 8435 39423
rect 8677 39389 8711 39423
rect 11621 39389 11655 39423
rect 12173 39389 12207 39423
rect 12449 39389 12483 39423
rect 14565 39389 14599 39423
rect 15853 39389 15887 39423
rect 16957 39389 16991 39423
rect 17785 39389 17819 39423
rect 18153 39389 18187 39423
rect 21833 39389 21867 39423
rect 24225 39389 24259 39423
rect 26985 39389 27019 39423
rect 28181 39389 28215 39423
rect 28273 39389 28307 39423
rect 28549 39389 28583 39423
rect 30849 39389 30883 39423
rect 31033 39389 31067 39423
rect 34897 39389 34931 39423
rect 36185 39389 36219 39423
rect 37197 39389 37231 39423
rect 37289 39389 37323 39423
rect 40785 39389 40819 39423
rect 41613 39389 41647 39423
rect 41981 39389 42015 39423
rect 43361 39389 43395 39423
rect 45201 39389 45235 39423
rect 47501 39389 47535 39423
rect 47685 39389 47719 39423
rect 49893 39389 49927 39423
rect 50169 39389 50203 39423
rect 50445 39389 50479 39423
rect 51641 39389 51675 39423
rect 54493 39389 54527 39423
rect 54585 39389 54619 39423
rect 55413 39389 55447 39423
rect 56241 39389 56275 39423
rect 57161 39389 57195 39423
rect 57345 39389 57379 39423
rect 59369 39389 59403 39423
rect 60013 39389 60047 39423
rect 30297 39321 30331 39355
rect 47041 39321 47075 39355
rect 51089 39321 51123 39355
rect 7849 39253 7883 39287
rect 10977 39253 11011 39287
rect 13921 39253 13955 39287
rect 14013 39253 14047 39287
rect 17141 39253 17175 39287
rect 21281 39253 21315 39287
rect 33701 39253 33735 39287
rect 35449 39253 35483 39287
rect 40233 39253 40267 39287
rect 41061 39253 41095 39287
rect 42625 39253 42659 39287
rect 44833 39253 44867 39287
rect 54033 39253 54067 39287
rect 56517 39253 56551 39287
rect 8217 39049 8251 39083
rect 12633 39049 12667 39083
rect 18705 39049 18739 39083
rect 19441 39049 19475 39083
rect 29272 39049 29306 39083
rect 43545 39049 43579 39083
rect 45845 39049 45879 39083
rect 47685 39049 47719 39083
rect 50445 39049 50479 39083
rect 54217 39049 54251 39083
rect 54769 39049 54803 39083
rect 57332 39049 57366 39083
rect 58817 39049 58851 39083
rect 58909 39049 58943 39083
rect 24685 38981 24719 39015
rect 26893 38981 26927 39015
rect 31677 38981 31711 39015
rect 32413 38981 32447 39015
rect 34161 38981 34195 39015
rect 39313 38981 39347 39015
rect 55597 38981 55631 39015
rect 6469 38913 6503 38947
rect 9413 38913 9447 38947
rect 10333 38913 10367 38947
rect 13093 38913 13127 38947
rect 13185 38913 13219 38947
rect 14473 38913 14507 38947
rect 15301 38913 15335 38947
rect 15393 38913 15427 38947
rect 16221 38913 16255 38947
rect 19901 38913 19935 38947
rect 19993 38913 20027 38947
rect 20729 38913 20763 38947
rect 20821 38913 20855 38947
rect 21649 38913 21683 38947
rect 24501 38913 24535 38947
rect 25145 38913 25179 38947
rect 25329 38913 25363 38947
rect 29009 38913 29043 38947
rect 30757 38913 30791 38947
rect 31493 38913 31527 38947
rect 33057 38913 33091 38947
rect 35909 38913 35943 38947
rect 37289 38913 37323 38947
rect 37381 38913 37415 38947
rect 38301 38913 38335 38947
rect 39037 38913 39071 38947
rect 39957 38913 39991 38947
rect 40601 38913 40635 38947
rect 40693 38913 40727 38947
rect 42993 38913 43027 38947
rect 44097 38913 44131 38947
rect 45201 38913 45235 38947
rect 45937 38913 45971 38947
rect 48329 38913 48363 38947
rect 49157 38913 49191 38947
rect 49341 38913 49375 38947
rect 50905 38913 50939 38947
rect 50997 38913 51031 38947
rect 52469 38913 52503 38947
rect 55229 38913 55263 38947
rect 55413 38913 55447 38947
rect 56333 38913 56367 38947
rect 57069 38913 57103 38947
rect 59461 38913 59495 38947
rect 10057 38845 10091 38879
rect 14289 38845 14323 38879
rect 19349 38845 19383 38879
rect 19809 38845 19843 38879
rect 21465 38845 21499 38879
rect 22477 38845 22511 38879
rect 23581 38845 23615 38879
rect 24225 38845 24259 38879
rect 25053 38845 25087 38879
rect 25513 38845 25547 38879
rect 26157 38845 26191 38879
rect 26341 38845 26375 38879
rect 32321 38845 32355 38879
rect 32873 38845 32907 38879
rect 38025 38845 38059 38879
rect 39773 38845 39807 38879
rect 40509 38845 40543 38879
rect 43269 38845 43303 38879
rect 49065 38845 49099 38879
rect 50261 38845 50295 38879
rect 52285 38845 52319 38879
rect 56149 38845 56183 38879
rect 59277 38845 59311 38879
rect 6745 38777 6779 38811
rect 9229 38777 9263 38811
rect 12081 38777 12115 38811
rect 13001 38777 13035 38811
rect 15669 38777 15703 38811
rect 16773 38777 16807 38811
rect 18521 38777 18555 38811
rect 20637 38777 20671 38811
rect 21925 38777 21959 38811
rect 24317 38777 24351 38811
rect 32781 38777 32815 38811
rect 35633 38777 35667 38811
rect 37197 38777 37231 38811
rect 38485 38777 38519 38811
rect 43913 38777 43947 38811
rect 45477 38777 45511 38811
rect 46213 38777 46247 38811
rect 50813 38777 50847 38811
rect 52745 38777 52779 38811
rect 8861 38709 8895 38743
rect 9321 38709 9355 38743
rect 13921 38709 13955 38743
rect 14381 38709 14415 38743
rect 14841 38709 14875 38743
rect 15209 38709 15243 38743
rect 20269 38709 20303 38743
rect 21097 38709 21131 38743
rect 21557 38709 21591 38743
rect 23029 38709 23063 38743
rect 23857 38709 23891 38743
rect 30849 38709 30883 38743
rect 31217 38709 31251 38743
rect 31309 38709 31343 38743
rect 36829 38709 36863 38743
rect 37657 38709 37691 38743
rect 38117 38709 38151 38743
rect 39681 38709 39715 38743
rect 40141 38709 40175 38743
rect 41521 38709 41555 38743
rect 44005 38709 44039 38743
rect 45385 38709 45419 38743
rect 47777 38709 47811 38743
rect 48697 38709 48731 38743
rect 51733 38709 51767 38743
rect 55137 38709 55171 38743
rect 55781 38709 55815 38743
rect 56241 38709 56275 38743
rect 59369 38709 59403 38743
rect 6929 38505 6963 38539
rect 7297 38505 7331 38539
rect 8125 38505 8159 38539
rect 10977 38505 11011 38539
rect 11713 38505 11747 38539
rect 15301 38505 15335 38539
rect 16497 38505 16531 38539
rect 21097 38505 21131 38539
rect 23305 38505 23339 38539
rect 25145 38505 25179 38539
rect 35449 38505 35483 38539
rect 35817 38505 35851 38539
rect 38485 38505 38519 38539
rect 41889 38505 41923 38539
rect 42349 38505 42383 38539
rect 45385 38505 45419 38539
rect 46121 38505 46155 38539
rect 46489 38505 46523 38539
rect 50445 38505 50479 38539
rect 50997 38505 51031 38539
rect 23673 38437 23707 38471
rect 29929 38437 29963 38471
rect 35909 38437 35943 38471
rect 37013 38437 37047 38471
rect 39589 38437 39623 38471
rect 48973 38437 49007 38471
rect 55505 38437 55539 38471
rect 8585 38369 8619 38403
rect 10609 38369 10643 38403
rect 12081 38369 12115 38403
rect 12909 38369 12943 38403
rect 13369 38369 13403 38403
rect 17233 38369 17267 38403
rect 17417 38369 17451 38403
rect 21557 38369 21591 38403
rect 26801 38369 26835 38403
rect 27261 38369 27295 38403
rect 29285 38369 29319 38403
rect 30481 38369 30515 38403
rect 31033 38369 31067 38403
rect 31585 38369 31619 38403
rect 33241 38369 33275 38403
rect 36461 38369 36495 38403
rect 36737 38369 36771 38403
rect 39313 38369 39347 38403
rect 42257 38369 42291 38403
rect 42717 38369 42751 38403
rect 43269 38369 43303 38403
rect 45293 38369 45327 38403
rect 48697 38369 48731 38403
rect 7389 38301 7423 38335
rect 7573 38301 7607 38335
rect 7941 38301 7975 38335
rect 8033 38301 8067 38335
rect 8861 38301 8895 38335
rect 11529 38301 11563 38335
rect 12173 38301 12207 38335
rect 12265 38301 12299 38335
rect 12633 38301 12667 38335
rect 12817 38301 12851 38335
rect 13645 38301 13679 38335
rect 15853 38301 15887 38335
rect 16589 38301 16623 38335
rect 16681 38301 16715 38335
rect 17693 38301 17727 38335
rect 19349 38301 19383 38335
rect 19625 38301 19659 38335
rect 21833 38301 21867 38335
rect 23397 38301 23431 38335
rect 26893 38301 26927 38335
rect 26985 38301 27019 38335
rect 27813 38301 27847 38335
rect 29377 38301 29411 38335
rect 29469 38301 29503 38335
rect 31125 38301 31159 38335
rect 31309 38301 31343 38335
rect 33517 38301 33551 38335
rect 34989 38301 35023 38335
rect 35173 38301 35207 38335
rect 35357 38301 35391 38335
rect 42533 38301 42567 38335
rect 45017 38301 45051 38335
rect 45937 38301 45971 38335
rect 46581 38301 46615 38335
rect 46673 38301 46707 38335
rect 47041 38301 47075 38335
rect 51089 38301 51123 38335
rect 51181 38301 51215 38335
rect 52745 38301 52779 38335
rect 53113 38301 53147 38335
rect 54861 38301 54895 38335
rect 55137 38301 55171 38335
rect 55229 38301 55263 38335
rect 57805 38301 57839 38335
rect 58081 38301 58115 38335
rect 59829 38301 59863 38335
rect 8493 38233 8527 38267
rect 13277 38233 13311 38267
rect 28917 38233 28951 38267
rect 15117 38165 15151 38199
rect 16129 38165 16163 38199
rect 19165 38165 19199 38199
rect 26433 38165 26467 38199
rect 30665 38165 30699 38199
rect 32229 38165 32263 38199
rect 41061 38165 41095 38199
rect 43545 38165 43579 38199
rect 47685 38165 47719 38199
rect 50629 38165 50663 38199
rect 52193 38165 52227 38199
rect 56977 38165 57011 38199
rect 9597 37961 9631 37995
rect 10425 37961 10459 37995
rect 14289 37961 14323 37995
rect 15779 37961 15813 37995
rect 17233 37961 17267 37995
rect 24672 37961 24706 37995
rect 28089 37961 28123 37995
rect 44189 37961 44223 37995
rect 44465 37961 44499 37995
rect 46397 37961 46431 37995
rect 50156 37961 50190 37995
rect 51733 37961 51767 37995
rect 54401 37961 54435 37995
rect 55781 37961 55815 37995
rect 18705 37893 18739 37927
rect 22937 37893 22971 37927
rect 34253 37893 34287 37927
rect 38945 37893 38979 37927
rect 42165 37893 42199 37927
rect 6469 37825 6503 37859
rect 8217 37825 8251 37859
rect 9413 37825 9447 37859
rect 10241 37825 10275 37859
rect 10977 37825 11011 37859
rect 16037 37825 16071 37859
rect 19257 37825 19291 37859
rect 20545 37825 20579 37859
rect 23489 37825 23523 37859
rect 24409 37825 24443 37859
rect 26249 37825 26283 37859
rect 28641 37825 28675 37859
rect 29929 37825 29963 37859
rect 30113 37825 30147 37859
rect 32045 37825 32079 37859
rect 34897 37825 34931 37859
rect 37105 37825 37139 37859
rect 37197 37825 37231 37859
rect 40417 37825 40451 37859
rect 43637 37825 43671 37859
rect 45017 37825 45051 37859
rect 48881 37825 48915 37859
rect 53757 37825 53791 37859
rect 55137 37825 55171 37859
rect 57897 37825 57931 37859
rect 59737 37825 59771 37859
rect 63693 37825 63727 37859
rect 63785 37825 63819 37859
rect 9137 37757 9171 37791
rect 16221 37757 16255 37791
rect 18521 37757 18555 37791
rect 19165 37757 19199 37791
rect 23305 37757 23339 37791
rect 32689 37757 32723 37791
rect 35357 37757 35391 37791
rect 43729 37757 43763 37791
rect 44833 37757 44867 37791
rect 48145 37757 48179 37791
rect 49893 37757 49927 37791
rect 53481 37757 53515 37791
rect 59921 37757 59955 37791
rect 6745 37689 6779 37723
rect 9229 37689 9263 37723
rect 10885 37689 10919 37723
rect 19073 37689 19107 37723
rect 20821 37689 20855 37723
rect 26525 37689 26559 37723
rect 28457 37689 28491 37723
rect 29837 37689 29871 37723
rect 31769 37689 31803 37723
rect 37473 37689 37507 37723
rect 40693 37689 40727 37723
rect 47869 37689 47903 37723
rect 53205 37689 53239 37723
rect 53941 37689 53975 37723
rect 54033 37689 54067 37723
rect 55321 37689 55355 37723
rect 55413 37689 55447 37723
rect 55873 37689 55907 37723
rect 57621 37689 57655 37723
rect 59461 37689 59495 37723
rect 63877 37689 63911 37723
rect 8769 37621 8803 37655
rect 9965 37621 9999 37655
rect 10057 37621 10091 37655
rect 10793 37621 10827 37655
rect 22293 37621 22327 37655
rect 23397 37621 23431 37655
rect 26157 37621 26191 37655
rect 27997 37621 28031 37655
rect 28549 37621 28583 37655
rect 29469 37621 29503 37655
rect 30297 37621 30331 37655
rect 32137 37621 32171 37655
rect 34621 37621 34655 37655
rect 34713 37621 34747 37655
rect 43821 37621 43855 37655
rect 44925 37621 44959 37655
rect 48237 37621 48271 37655
rect 48605 37621 48639 37655
rect 48697 37621 48731 37655
rect 51641 37621 51675 37655
rect 57989 37621 58023 37655
rect 60565 37621 60599 37655
rect 64245 37621 64279 37655
rect 18705 37417 18739 37451
rect 19073 37417 19107 37451
rect 21465 37417 21499 37451
rect 21833 37417 21867 37451
rect 23857 37417 23891 37451
rect 24225 37417 24259 37451
rect 26893 37417 26927 37451
rect 27261 37417 27295 37451
rect 31125 37417 31159 37451
rect 31585 37417 31619 37451
rect 31953 37417 31987 37451
rect 32045 37417 32079 37451
rect 34529 37417 34563 37451
rect 34897 37417 34931 37451
rect 35449 37417 35483 37451
rect 35817 37417 35851 37451
rect 39313 37417 39347 37451
rect 40417 37417 40451 37451
rect 40877 37417 40911 37451
rect 40969 37417 41003 37451
rect 41429 37417 41463 37451
rect 46213 37417 46247 37451
rect 46673 37417 46707 37451
rect 47501 37417 47535 37451
rect 47869 37417 47903 37451
rect 50169 37417 50203 37451
rect 50629 37417 50663 37451
rect 51089 37417 51123 37451
rect 51549 37417 51583 37451
rect 53021 37417 53055 37451
rect 53481 37417 53515 37451
rect 57345 37417 57379 37451
rect 57713 37417 57747 37451
rect 57805 37417 57839 37451
rect 58173 37417 58207 37451
rect 58541 37417 58575 37451
rect 58633 37417 58667 37451
rect 59369 37417 59403 37451
rect 59737 37417 59771 37451
rect 59921 37417 59955 37451
rect 60289 37417 60323 37451
rect 64889 37417 64923 37451
rect 8769 37349 8803 37383
rect 19165 37349 19199 37383
rect 21925 37349 21959 37383
rect 29653 37349 29687 37383
rect 36737 37349 36771 37383
rect 40509 37349 40543 37383
rect 47409 37349 47443 37383
rect 51641 37349 51675 37383
rect 53389 37349 53423 37383
rect 8493 37281 8527 37315
rect 10517 37281 10551 37315
rect 13553 37281 13587 37315
rect 16589 37281 16623 37315
rect 24317 37281 24351 37315
rect 27353 37281 27387 37315
rect 27721 37281 27755 37315
rect 28365 37281 28399 37315
rect 29377 37281 29411 37315
rect 34989 37281 35023 37315
rect 39681 37281 39715 37315
rect 41337 37281 41371 37315
rect 46305 37281 46339 37315
rect 50721 37281 50755 37315
rect 54493 37281 54527 37315
rect 54953 37281 54987 37315
rect 59277 37281 59311 37315
rect 60381 37281 60415 37315
rect 63141 37281 63175 37315
rect 65625 37281 65659 37315
rect 13829 37213 13863 37247
rect 15301 37213 15335 37247
rect 16865 37213 16899 37247
rect 18337 37213 18371 37247
rect 19257 37213 19291 37247
rect 22017 37213 22051 37247
rect 24501 37213 24535 37247
rect 27445 37213 27479 37247
rect 32137 37213 32171 37247
rect 34253 37213 34287 37247
rect 34437 37213 34471 37247
rect 35909 37213 35943 37247
rect 36093 37213 36127 37247
rect 38485 37213 38519 37247
rect 39773 37213 39807 37247
rect 39865 37213 39899 37247
rect 40325 37213 40359 37247
rect 41521 37213 41555 37247
rect 46121 37213 46155 37247
rect 47317 37213 47351 37247
rect 50537 37213 50571 37247
rect 51457 37213 51491 37247
rect 52929 37213 52963 37247
rect 53573 37213 53607 37247
rect 57897 37213 57931 37247
rect 58725 37213 58759 37247
rect 59093 37213 59127 37247
rect 60473 37213 60507 37247
rect 63417 37213 63451 37247
rect 35357 37145 35391 37179
rect 52009 37145 52043 37179
rect 56425 37077 56459 37111
rect 65073 37077 65107 37111
rect 63877 36873 63911 36907
rect 64337 36737 64371 36771
rect 64429 36737 64463 36771
rect 65993 36737 66027 36771
rect 64245 36601 64279 36635
rect 65441 36533 65475 36567
rect 65625 36329 65659 36363
rect 63877 36125 63911 36159
rect 64153 36125 64187 36159
rect 64705 35785 64739 35819
rect 63969 35649 64003 35683
rect 64153 35649 64187 35683
rect 65349 35649 65383 35683
rect 64245 35581 64279 35615
rect 65073 35581 65107 35615
rect 65165 35513 65199 35547
rect 64613 35445 64647 35479
rect 65625 34697 65659 34731
rect 63877 34493 63911 34527
rect 64153 34425 64187 34459
rect 63969 34153 64003 34187
rect 64337 34017 64371 34051
rect 65073 34017 65107 34051
rect 65625 34017 65659 34051
rect 64429 33949 64463 33983
rect 64613 33949 64647 33983
rect 64705 33473 64739 33507
rect 64981 33405 65015 33439
rect 65993 33405 66027 33439
rect 64889 33337 64923 33371
rect 65349 33269 65383 33303
rect 65441 33269 65475 33303
rect 63969 32861 64003 32895
rect 64245 32861 64279 32895
rect 65717 32725 65751 32759
rect 64705 32521 64739 32555
rect 64981 32521 65015 32555
rect 64153 32385 64187 32419
rect 65441 32385 65475 32419
rect 65533 32385 65567 32419
rect 64245 32317 64279 32351
rect 65349 32317 65383 32351
rect 64337 32249 64371 32283
rect 64797 32249 64831 32283
rect 65441 31977 65475 32011
rect 64153 31909 64187 31943
rect 64061 31841 64095 31875
rect 64613 31365 64647 31399
rect 65257 31297 65291 31331
rect 65073 31229 65107 31263
rect 64981 31161 65015 31195
rect 64061 30753 64095 30787
rect 64337 30685 64371 30719
rect 65809 30549 65843 30583
rect 64613 30345 64647 30379
rect 65073 30209 65107 30243
rect 65257 30209 65291 30243
rect 65993 30141 66027 30175
rect 64981 30073 65015 30107
rect 65441 30073 65475 30107
rect 64981 29733 65015 29767
rect 64889 29665 64923 29699
rect 65441 29665 65475 29699
rect 65165 29597 65199 29631
rect 65993 29597 66027 29631
rect 64521 29461 64555 29495
rect 64061 29121 64095 29155
rect 64337 29121 64371 29155
rect 65809 29121 65843 29155
rect 65073 28713 65107 28747
rect 64705 28645 64739 28679
rect 64613 28577 64647 28611
rect 64521 28509 64555 28543
rect 64613 27013 64647 27047
rect 65165 26945 65199 26979
rect 65073 26877 65107 26911
rect 64981 26809 65015 26843
rect 64061 26333 64095 26367
rect 64337 26333 64371 26367
rect 65809 26197 65843 26231
rect 64613 25993 64647 26027
rect 65073 25857 65107 25891
rect 65257 25857 65291 25891
rect 65993 25789 66027 25823
rect 64981 25653 65015 25687
rect 65441 25653 65475 25687
rect 64337 25313 64371 25347
rect 64981 25313 65015 25347
rect 65441 25313 65475 25347
rect 65073 25245 65107 25279
rect 65165 25245 65199 25279
rect 65993 25245 66027 25279
rect 64613 25109 64647 25143
rect 63877 24701 63911 24735
rect 65165 24565 65199 24599
rect 64337 24293 64371 24327
rect 64061 24157 64095 24191
rect 65809 24021 65843 24055
rect 63877 23613 63911 23647
rect 65165 23477 65199 23511
rect 65257 23273 65291 23307
rect 64797 23205 64831 23239
rect 64061 23137 64095 23171
rect 64889 23137 64923 23171
rect 64705 23069 64739 23103
rect 64613 22729 64647 22763
rect 65809 22185 65843 22219
rect 64061 21981 64095 22015
rect 64337 21981 64371 22015
rect 66085 21505 66119 21539
rect 65073 21437 65107 21471
rect 64797 21301 64831 21335
rect 65441 21301 65475 21335
rect 64613 21097 64647 21131
rect 64981 21097 65015 21131
rect 65073 21029 65107 21063
rect 65533 21029 65567 21063
rect 65257 20893 65291 20927
rect 65809 20757 65843 20791
rect 64613 20485 64647 20519
rect 65257 20417 65291 20451
rect 65073 20349 65107 20383
rect 64981 20213 65015 20247
rect 64061 19873 64095 19907
rect 64337 19805 64371 19839
rect 65809 19669 65843 19703
rect 64613 19465 64647 19499
rect 65257 19329 65291 19363
rect 65073 19261 65107 19295
rect 65993 19261 66027 19295
rect 64981 19193 65015 19227
rect 65441 19193 65475 19227
rect 64981 18785 65015 18819
rect 65441 18785 65475 18819
rect 65073 18717 65107 18751
rect 65257 18717 65291 18751
rect 65993 18717 66027 18751
rect 64613 18581 64647 18615
rect 64061 18241 64095 18275
rect 64337 18241 64371 18275
rect 65809 18037 65843 18071
rect 64889 17833 64923 17867
rect 65349 17833 65383 17867
rect 65717 17833 65751 17867
rect 64797 17765 64831 17799
rect 64705 17629 64739 17663
rect 65809 17629 65843 17663
rect 65901 17629 65935 17663
rect 65257 17561 65291 17595
rect 64521 17289 64555 17323
rect 65441 16609 65475 16643
rect 66085 16405 66119 16439
rect 65349 16133 65383 16167
rect 64705 16065 64739 16099
rect 65901 16065 65935 16099
rect 64889 15997 64923 16031
rect 65717 15997 65751 16031
rect 65809 15929 65843 15963
rect 64797 15861 64831 15895
rect 65257 15861 65291 15895
rect 64613 15657 64647 15691
rect 64337 14977 64371 15011
rect 64061 14909 64095 14943
rect 65809 14773 65843 14807
rect 65809 13481 65843 13515
rect 64337 13413 64371 13447
rect 64061 13277 64095 13311
rect 65993 12801 66027 12835
rect 65441 12597 65475 12631
rect 64061 12189 64095 12223
rect 64337 12189 64371 12223
rect 66085 12189 66119 12223
rect 64613 11849 64647 11883
rect 65165 11713 65199 11747
rect 64981 11645 65015 11679
rect 65073 11509 65107 11543
rect 64521 11305 64555 11339
rect 64889 11237 64923 11271
rect 64981 11169 65015 11203
rect 65165 11101 65199 11135
rect 65165 10625 65199 10659
rect 65073 10557 65107 10591
rect 64613 10421 64647 10455
rect 64981 10421 65015 10455
rect 64981 10217 65015 10251
rect 64797 10013 64831 10047
rect 64889 10013 64923 10047
rect 65349 9877 65383 9911
rect 65993 9469 66027 9503
rect 65441 9333 65475 9367
rect 64061 8925 64095 8959
rect 64337 8925 64371 8959
rect 65809 8789 65843 8823
rect 64613 8585 64647 8619
rect 65257 8449 65291 8483
rect 65993 8449 66027 8483
rect 65073 8381 65107 8415
rect 64981 8313 65015 8347
rect 65441 8313 65475 8347
rect 65809 8041 65843 8075
rect 64061 7905 64095 7939
rect 64337 7837 64371 7871
rect 64429 7497 64463 7531
rect 64613 7497 64647 7531
rect 65073 7361 65107 7395
rect 65257 7361 65291 7395
rect 64981 7293 65015 7327
rect 65993 7293 66027 7327
rect 65441 7157 65475 7191
rect 64797 6953 64831 6987
rect 65625 6953 65659 6987
rect 63877 6817 63911 6851
rect 64705 6817 64739 6851
rect 65717 6817 65751 6851
rect 64153 6749 64187 6783
rect 64613 6749 64647 6783
rect 65809 6749 65843 6783
rect 65165 6681 65199 6715
rect 65257 6613 65291 6647
rect 64429 6409 64463 6443
rect 64705 6341 64739 6375
rect 65257 6273 65291 6307
rect 65165 6205 65199 6239
rect 65073 6069 65107 6103
rect 64153 5865 64187 5899
rect 64705 5865 64739 5899
rect 64245 5797 64279 5831
rect 65257 5729 65291 5763
rect 64061 5661 64095 5695
rect 65349 5661 65383 5695
rect 65441 5661 65475 5695
rect 64613 5593 64647 5627
rect 64889 5525 64923 5559
rect 63877 5185 63911 5219
rect 64153 5185 64187 5219
rect 65625 4981 65659 5015
rect 65809 4777 65843 4811
rect 64337 4709 64371 4743
rect 64061 4641 64095 4675
rect 63877 4029 63911 4063
rect 64153 3961 64187 3995
rect 65625 3893 65659 3927
rect 64705 3689 64739 3723
rect 64245 3621 64279 3655
rect 65073 3621 65107 3655
rect 63969 3485 64003 3519
rect 64153 3485 64187 3519
rect 65165 3485 65199 3519
rect 65349 3485 65383 3519
rect 64613 3417 64647 3451
rect 63969 3145 64003 3179
rect 64061 3009 64095 3043
rect 65809 3009 65843 3043
rect 64337 2873 64371 2907
rect 64613 2601 64647 2635
rect 65165 2601 65199 2635
rect 65073 2533 65107 2567
rect 64245 2465 64279 2499
rect 64061 2397 64095 2431
rect 64153 2397 64187 2431
rect 65257 2397 65291 2431
rect 64705 2329 64739 2363
rect 65441 2057 65475 2091
rect 64613 1989 64647 2023
rect 65257 1921 65291 1955
rect 65993 1921 66027 1955
rect 64981 1853 65015 1887
rect 65073 1853 65107 1887
rect 65441 1513 65475 1547
rect 64705 1309 64739 1343
rect 65993 1309 66027 1343
rect 65441 969 65475 1003
rect 65993 833 66027 867
<< metal1 >>
rect 27706 44820 27712 44872
rect 27764 44860 27770 44872
rect 28810 44860 28816 44872
rect 27764 44832 28816 44860
rect 27764 44820 27770 44832
rect 28810 44820 28816 44832
rect 28868 44860 28874 44872
rect 30926 44860 30932 44872
rect 28868 44832 30932 44860
rect 28868 44820 28874 44832
rect 30926 44820 30932 44832
rect 30984 44820 30990 44872
rect 16758 44752 16764 44804
rect 16816 44792 16822 44804
rect 21726 44792 21732 44804
rect 16816 44764 21732 44792
rect 16816 44752 16822 44764
rect 21726 44752 21732 44764
rect 21784 44752 21790 44804
rect 24854 44752 24860 44804
rect 24912 44792 24918 44804
rect 33502 44792 33508 44804
rect 24912 44764 33508 44792
rect 24912 44752 24918 44764
rect 33502 44752 33508 44764
rect 33560 44752 33566 44804
rect 17310 44684 17316 44736
rect 17368 44724 17374 44736
rect 24026 44724 24032 44736
rect 17368 44696 24032 44724
rect 17368 44684 17374 44696
rect 24026 44684 24032 44696
rect 24084 44684 24090 44736
rect 29178 44684 29184 44736
rect 29236 44724 29242 44736
rect 40402 44724 40408 44736
rect 29236 44696 40408 44724
rect 29236 44684 29242 44696
rect 40402 44684 40408 44696
rect 40460 44684 40466 44736
rect 552 44634 66424 44656
rect 552 44582 1998 44634
rect 2050 44582 2062 44634
rect 2114 44582 2126 44634
rect 2178 44582 2190 44634
rect 2242 44582 2254 44634
rect 2306 44582 50998 44634
rect 51050 44582 51062 44634
rect 51114 44582 51126 44634
rect 51178 44582 51190 44634
rect 51242 44582 51254 44634
rect 51306 44582 66424 44634
rect 552 44560 66424 44582
rect 6178 44480 6184 44532
rect 6236 44480 6242 44532
rect 6730 44480 6736 44532
rect 6788 44480 6794 44532
rect 7282 44480 7288 44532
rect 7340 44480 7346 44532
rect 7834 44480 7840 44532
rect 7892 44480 7898 44532
rect 8386 44480 8392 44532
rect 8444 44480 8450 44532
rect 8938 44480 8944 44532
rect 8996 44480 9002 44532
rect 9490 44480 9496 44532
rect 9548 44480 9554 44532
rect 10042 44480 10048 44532
rect 10100 44480 10106 44532
rect 10594 44480 10600 44532
rect 10652 44480 10658 44532
rect 12250 44480 12256 44532
rect 12308 44480 12314 44532
rect 12526 44480 12532 44532
rect 12584 44480 12590 44532
rect 12802 44480 12808 44532
rect 12860 44480 12866 44532
rect 13538 44480 13544 44532
rect 13596 44480 13602 44532
rect 13814 44480 13820 44532
rect 13872 44480 13878 44532
rect 15470 44480 15476 44532
rect 15528 44480 15534 44532
rect 15930 44480 15936 44532
rect 15988 44480 15994 44532
rect 16206 44480 16212 44532
rect 16264 44480 16270 44532
rect 16666 44480 16672 44532
rect 16724 44480 16730 44532
rect 16942 44480 16948 44532
rect 17000 44480 17006 44532
rect 17218 44480 17224 44532
rect 17276 44480 17282 44532
rect 20070 44520 20076 44532
rect 19306 44492 20076 44520
rect 19306 44452 19334 44492
rect 20070 44480 20076 44492
rect 20128 44480 20134 44532
rect 21726 44480 21732 44532
rect 21784 44520 21790 44532
rect 30837 44523 30895 44529
rect 30837 44520 30849 44523
rect 21784 44492 30849 44520
rect 21784 44480 21790 44492
rect 30837 44489 30849 44492
rect 30883 44489 30895 44523
rect 30837 44483 30895 44489
rect 17788 44424 19334 44452
rect 24949 44455 25007 44461
rect 10965 44319 11023 44325
rect 10965 44285 10977 44319
rect 11011 44316 11023 44319
rect 12250 44316 12256 44328
rect 11011 44288 12256 44316
rect 11011 44285 11023 44288
rect 10965 44279 11023 44285
rect 12250 44276 12256 44288
rect 12308 44276 12314 44328
rect 14366 44276 14372 44328
rect 14424 44316 14430 44328
rect 14645 44319 14703 44325
rect 14645 44316 14657 44319
rect 14424 44288 14657 44316
rect 14424 44276 14430 44288
rect 14645 44285 14657 44288
rect 14691 44285 14703 44319
rect 14645 44279 14703 44285
rect 17699 44319 17757 44325
rect 17699 44285 17711 44319
rect 17745 44316 17757 44319
rect 17788 44316 17816 44424
rect 24949 44421 24961 44455
rect 24995 44452 25007 44455
rect 26418 44452 26424 44464
rect 24995 44424 26424 44452
rect 24995 44421 25007 44424
rect 24949 44415 25007 44421
rect 26418 44412 26424 44424
rect 26476 44412 26482 44464
rect 30377 44455 30435 44461
rect 30377 44452 30389 44455
rect 27448 44424 30389 44452
rect 17862 44344 17868 44396
rect 17920 44384 17926 44396
rect 19337 44387 19395 44393
rect 19337 44384 19349 44387
rect 17920 44356 18644 44384
rect 17920 44344 17926 44356
rect 17745 44288 17816 44316
rect 17745 44285 17757 44288
rect 17699 44279 17757 44285
rect 18506 44276 18512 44328
rect 18564 44276 18570 44328
rect 18616 44316 18644 44356
rect 19076 44356 19349 44384
rect 19076 44316 19104 44356
rect 19337 44353 19349 44356
rect 19383 44384 19395 44387
rect 20533 44387 20591 44393
rect 19383 44356 20208 44384
rect 19383 44353 19395 44356
rect 19337 44347 19395 44353
rect 18616 44288 19104 44316
rect 19150 44276 19156 44328
rect 19208 44316 19214 44328
rect 20073 44319 20131 44325
rect 20073 44316 20085 44319
rect 19208 44288 20085 44316
rect 19208 44276 19214 44288
rect 20073 44285 20085 44288
rect 20119 44285 20131 44319
rect 20073 44279 20131 44285
rect 10594 44208 10600 44260
rect 10652 44248 10658 44260
rect 11701 44251 11759 44257
rect 11701 44248 11713 44251
rect 10652 44220 11713 44248
rect 10652 44208 10658 44220
rect 11701 44217 11713 44220
rect 11747 44217 11759 44251
rect 11701 44211 11759 44217
rect 12069 44251 12127 44257
rect 12069 44217 12081 44251
rect 12115 44217 12127 44251
rect 14182 44248 14188 44260
rect 12069 44211 12127 44217
rect 12406 44220 14188 44248
rect 11606 44140 11612 44192
rect 11664 44140 11670 44192
rect 12084 44180 12112 44211
rect 12406 44180 12434 44220
rect 14182 44208 14188 44220
rect 14240 44208 14246 44260
rect 14461 44251 14519 44257
rect 14461 44217 14473 44251
rect 14507 44248 14519 44251
rect 18874 44248 18880 44260
rect 14507 44220 18880 44248
rect 14507 44217 14519 44220
rect 14461 44211 14519 44217
rect 18874 44208 18880 44220
rect 18932 44208 18938 44260
rect 19061 44251 19119 44257
rect 19061 44217 19073 44251
rect 19107 44248 19119 44251
rect 19521 44251 19579 44257
rect 19521 44248 19533 44251
rect 19107 44220 19533 44248
rect 19107 44217 19119 44220
rect 19061 44211 19119 44217
rect 19521 44217 19533 44220
rect 19567 44217 19579 44251
rect 20180 44248 20208 44356
rect 20533 44353 20545 44387
rect 20579 44384 20591 44387
rect 22278 44384 22284 44396
rect 20579 44356 22284 44384
rect 20579 44353 20591 44356
rect 20533 44347 20591 44353
rect 22278 44344 22284 44356
rect 22336 44344 22342 44396
rect 22465 44387 22523 44393
rect 22465 44353 22477 44387
rect 22511 44384 22523 44387
rect 23934 44384 23940 44396
rect 22511 44356 23940 44384
rect 22511 44353 22523 44356
rect 22465 44347 22523 44353
rect 21085 44319 21143 44325
rect 21085 44285 21097 44319
rect 21131 44316 21143 44319
rect 22189 44319 22247 44325
rect 22189 44316 22201 44319
rect 21131 44288 22201 44316
rect 21131 44285 21143 44288
rect 21085 44279 21143 44285
rect 22189 44285 22201 44288
rect 22235 44285 22247 44319
rect 22189 44279 22247 44285
rect 20714 44248 20720 44260
rect 20180 44220 20720 44248
rect 19521 44211 19579 44217
rect 20714 44208 20720 44220
rect 20772 44248 20778 44260
rect 20990 44248 20996 44260
rect 20772 44220 20996 44248
rect 20772 44208 20778 44220
rect 20990 44208 20996 44220
rect 21048 44248 21054 44260
rect 21269 44251 21327 44257
rect 21269 44248 21281 44251
rect 21048 44220 21281 44248
rect 21048 44208 21054 44220
rect 21269 44217 21281 44220
rect 21315 44217 21327 44251
rect 21269 44211 21327 44217
rect 21450 44208 21456 44260
rect 21508 44248 21514 44260
rect 21637 44251 21695 44257
rect 21637 44248 21649 44251
rect 21508 44220 21649 44248
rect 21508 44208 21514 44220
rect 21637 44217 21649 44220
rect 21683 44248 21695 44251
rect 22480 44248 22508 44347
rect 23934 44344 23940 44356
rect 23992 44344 23998 44396
rect 25685 44387 25743 44393
rect 25685 44353 25697 44387
rect 25731 44384 25743 44387
rect 25731 44356 26740 44384
rect 25731 44353 25743 44356
rect 25685 44347 25743 44353
rect 22554 44276 22560 44328
rect 22612 44316 22618 44328
rect 23477 44319 23535 44325
rect 23477 44316 23489 44319
rect 22612 44288 23489 44316
rect 22612 44276 22618 44288
rect 23477 44285 23489 44288
rect 23523 44285 23535 44319
rect 23477 44279 23535 44285
rect 24026 44276 24032 44328
rect 24084 44276 24090 44328
rect 24397 44319 24455 44325
rect 24397 44285 24409 44319
rect 24443 44316 24455 44319
rect 26234 44316 26240 44328
rect 24443 44288 26240 44316
rect 24443 44285 24455 44288
rect 24397 44279 24455 44285
rect 26234 44276 26240 44288
rect 26292 44276 26298 44328
rect 26602 44276 26608 44328
rect 26660 44276 26666 44328
rect 26712 44316 26740 44356
rect 26786 44344 26792 44396
rect 26844 44344 26850 44396
rect 27448 44328 27476 44424
rect 30377 44421 30389 44424
rect 30423 44421 30435 44455
rect 30377 44415 30435 44421
rect 27522 44344 27528 44396
rect 27580 44344 27586 44396
rect 28813 44387 28871 44393
rect 28813 44353 28825 44387
rect 28859 44384 28871 44387
rect 28859 44356 30788 44384
rect 28859 44353 28871 44356
rect 28813 44347 28871 44353
rect 27430 44316 27436 44328
rect 26712 44288 27436 44316
rect 27430 44276 27436 44288
rect 27488 44276 27494 44328
rect 28261 44319 28319 44325
rect 28261 44285 28273 44319
rect 28307 44316 28319 44319
rect 28626 44316 28632 44328
rect 28307 44288 28632 44316
rect 28307 44285 28319 44288
rect 28261 44279 28319 44285
rect 28626 44276 28632 44288
rect 28684 44276 28690 44328
rect 30009 44319 30067 44325
rect 30009 44285 30021 44319
rect 30055 44316 30067 44319
rect 30466 44316 30472 44328
rect 30055 44288 30472 44316
rect 30055 44285 30067 44288
rect 30009 44279 30067 44285
rect 30466 44276 30472 44288
rect 30524 44276 30530 44328
rect 30760 44325 30788 44356
rect 30745 44319 30803 44325
rect 30745 44285 30757 44319
rect 30791 44285 30803 44319
rect 30852 44316 30880 44483
rect 30926 44480 30932 44532
rect 30984 44520 30990 44532
rect 30984 44492 35894 44520
rect 30984 44480 30990 44492
rect 35866 44452 35894 44492
rect 36538 44480 36544 44532
rect 36596 44520 36602 44532
rect 40221 44523 40279 44529
rect 36596 44492 38240 44520
rect 36596 44480 36602 44492
rect 38102 44452 38108 44464
rect 35866 44424 36952 44452
rect 33042 44344 33048 44396
rect 33100 44384 33106 44396
rect 33505 44387 33563 44393
rect 33505 44384 33517 44387
rect 33100 44356 33517 44384
rect 33100 44344 33106 44356
rect 33505 44353 33517 44356
rect 33551 44384 33563 44387
rect 34977 44387 35035 44393
rect 34977 44384 34989 44387
rect 33551 44356 34989 44384
rect 33551 44353 33563 44356
rect 33505 44347 33563 44353
rect 34977 44353 34989 44356
rect 35023 44384 35035 44387
rect 35710 44384 35716 44396
rect 35023 44356 35716 44384
rect 35023 44353 35035 44356
rect 34977 44347 35035 44353
rect 35710 44344 35716 44356
rect 35768 44344 35774 44396
rect 31297 44319 31355 44325
rect 31297 44316 31309 44319
rect 30852 44288 31309 44316
rect 30745 44279 30803 44285
rect 31297 44285 31309 44288
rect 31343 44316 31355 44319
rect 31846 44316 31852 44328
rect 31343 44288 31852 44316
rect 31343 44285 31355 44288
rect 31297 44279 31355 44285
rect 31846 44276 31852 44288
rect 31904 44316 31910 44328
rect 34238 44316 34244 44328
rect 31904 44288 34244 44316
rect 31904 44276 31910 44288
rect 34238 44276 34244 44288
rect 34296 44276 34302 44328
rect 35434 44276 35440 44328
rect 35492 44316 35498 44328
rect 36924 44325 36952 44424
rect 37200 44424 38108 44452
rect 37200 44393 37228 44424
rect 38102 44412 38108 44424
rect 38160 44412 38166 44464
rect 37185 44387 37243 44393
rect 37185 44353 37197 44387
rect 37231 44353 37243 44387
rect 37918 44384 37924 44396
rect 37185 44347 37243 44353
rect 37844 44356 37924 44384
rect 37844 44325 37872 44356
rect 37918 44344 37924 44356
rect 37976 44344 37982 44396
rect 38010 44344 38016 44396
rect 38068 44344 38074 44396
rect 38212 44384 38240 44492
rect 40221 44489 40233 44523
rect 40267 44520 40279 44523
rect 41598 44520 41604 44532
rect 40267 44492 41604 44520
rect 40267 44489 40279 44492
rect 40221 44483 40279 44489
rect 41598 44480 41604 44492
rect 41656 44520 41662 44532
rect 42518 44520 42524 44532
rect 41656 44492 42524 44520
rect 41656 44480 41662 44492
rect 42518 44480 42524 44492
rect 42576 44480 42582 44532
rect 38286 44412 38292 44464
rect 38344 44452 38350 44464
rect 39390 44452 39396 44464
rect 38344 44424 39396 44452
rect 38344 44412 38350 44424
rect 39390 44412 39396 44424
rect 39448 44452 39454 44464
rect 39448 44424 46428 44452
rect 39448 44412 39454 44424
rect 38212 44356 41000 44384
rect 35805 44319 35863 44325
rect 35805 44316 35817 44319
rect 35492 44288 35817 44316
rect 35492 44276 35498 44288
rect 35805 44285 35817 44288
rect 35851 44285 35863 44319
rect 35805 44279 35863 44285
rect 36909 44319 36967 44325
rect 36909 44285 36921 44319
rect 36955 44285 36967 44319
rect 36909 44279 36967 44285
rect 37829 44319 37887 44325
rect 37829 44285 37841 44319
rect 37875 44285 37887 44319
rect 37829 44279 37887 44285
rect 38286 44276 38292 44328
rect 38344 44276 38350 44328
rect 39669 44319 39727 44325
rect 39669 44285 39681 44319
rect 39715 44316 39727 44319
rect 39850 44316 39856 44328
rect 39715 44288 39856 44316
rect 39715 44285 39727 44288
rect 39669 44279 39727 44285
rect 39850 44276 39856 44288
rect 39908 44276 39914 44328
rect 40402 44276 40408 44328
rect 40460 44276 40466 44328
rect 40972 44325 41000 44356
rect 42518 44344 42524 44396
rect 42576 44384 42582 44396
rect 43070 44384 43076 44396
rect 42576 44356 43076 44384
rect 42576 44344 42582 44356
rect 43070 44344 43076 44356
rect 43128 44344 43134 44396
rect 43257 44387 43315 44393
rect 43257 44353 43269 44387
rect 43303 44384 43315 44387
rect 43990 44384 43996 44396
rect 43303 44356 43996 44384
rect 43303 44353 43315 44356
rect 43257 44347 43315 44353
rect 40957 44319 41015 44325
rect 40957 44285 40969 44319
rect 41003 44285 41015 44319
rect 43272 44316 43300 44347
rect 43990 44344 43996 44356
rect 44048 44344 44054 44396
rect 40957 44279 41015 44285
rect 41340 44288 43300 44316
rect 21683 44220 22508 44248
rect 21683 44217 21695 44220
rect 21637 44211 21695 44217
rect 23382 44208 23388 44260
rect 23440 44248 23446 44260
rect 23845 44251 23903 44257
rect 23845 44248 23857 44251
rect 23440 44220 23857 44248
rect 23440 44208 23446 44220
rect 23845 44217 23857 44220
rect 23891 44217 23903 44251
rect 24044 44248 24072 44276
rect 25869 44251 25927 44257
rect 25869 44248 25881 44251
rect 24044 44220 25881 44248
rect 23845 44211 23903 44217
rect 25869 44217 25881 44220
rect 25915 44217 25927 44251
rect 25869 44211 25927 44217
rect 26050 44208 26056 44260
rect 26108 44248 26114 44260
rect 26108 44220 29132 44248
rect 26108 44208 26114 44220
rect 12084 44152 12434 44180
rect 12526 44140 12532 44192
rect 12584 44180 12590 44192
rect 12894 44180 12900 44192
rect 12584 44152 12900 44180
rect 12584 44140 12590 44152
rect 12894 44140 12900 44152
rect 12952 44180 12958 44192
rect 14369 44183 14427 44189
rect 14369 44180 14381 44183
rect 12952 44152 14381 44180
rect 12952 44140 12958 44152
rect 14369 44149 14381 44152
rect 14415 44180 14427 44183
rect 14734 44180 14740 44192
rect 14415 44152 14740 44180
rect 14415 44149 14427 44152
rect 14369 44143 14427 44149
rect 14734 44140 14740 44152
rect 14792 44140 14798 44192
rect 14826 44140 14832 44192
rect 14884 44180 14890 44192
rect 15289 44183 15347 44189
rect 15289 44180 15301 44183
rect 14884 44152 15301 44180
rect 14884 44140 14890 44152
rect 15289 44149 15301 44152
rect 15335 44149 15347 44183
rect 15289 44143 15347 44149
rect 17405 44183 17463 44189
rect 17405 44149 17417 44183
rect 17451 44180 17463 44183
rect 17494 44180 17500 44192
rect 17451 44152 17500 44180
rect 17451 44149 17463 44152
rect 17405 44143 17463 44149
rect 17494 44140 17500 44152
rect 17552 44140 17558 44192
rect 17586 44140 17592 44192
rect 17644 44180 17650 44192
rect 17865 44183 17923 44189
rect 17865 44180 17877 44183
rect 17644 44152 17877 44180
rect 17644 44140 17650 44152
rect 17865 44149 17877 44152
rect 17911 44149 17923 44183
rect 17865 44143 17923 44149
rect 18693 44183 18751 44189
rect 18693 44149 18705 44183
rect 18739 44180 18751 44183
rect 18966 44180 18972 44192
rect 18739 44152 18972 44180
rect 18739 44149 18751 44152
rect 18693 44143 18751 44149
rect 18966 44140 18972 44152
rect 19024 44140 19030 44192
rect 19153 44183 19211 44189
rect 19153 44149 19165 44183
rect 19199 44180 19211 44183
rect 20254 44180 20260 44192
rect 19199 44152 20260 44180
rect 19199 44149 19211 44152
rect 19153 44143 19211 44149
rect 20254 44140 20260 44152
rect 20312 44140 20318 44192
rect 21542 44140 21548 44192
rect 21600 44180 21606 44192
rect 21821 44183 21879 44189
rect 21821 44180 21833 44183
rect 21600 44152 21833 44180
rect 21600 44140 21606 44152
rect 21821 44149 21833 44152
rect 21867 44149 21879 44183
rect 21821 44143 21879 44149
rect 22094 44140 22100 44192
rect 22152 44180 22158 44192
rect 22281 44183 22339 44189
rect 22281 44180 22293 44183
rect 22152 44152 22293 44180
rect 22152 44140 22158 44152
rect 22281 44149 22293 44152
rect 22327 44149 22339 44183
rect 22281 44143 22339 44149
rect 22462 44140 22468 44192
rect 22520 44180 22526 44192
rect 22925 44183 22983 44189
rect 22925 44180 22937 44183
rect 22520 44152 22937 44180
rect 22520 44140 22526 44152
rect 22925 44149 22937 44152
rect 22971 44149 22983 44183
rect 22925 44143 22983 44149
rect 25038 44140 25044 44192
rect 25096 44140 25102 44192
rect 25314 44140 25320 44192
rect 25372 44180 25378 44192
rect 25409 44183 25467 44189
rect 25409 44180 25421 44183
rect 25372 44152 25421 44180
rect 25372 44140 25378 44152
rect 25409 44149 25421 44152
rect 25455 44149 25467 44183
rect 25409 44143 25467 44149
rect 25498 44140 25504 44192
rect 25556 44140 25562 44192
rect 25590 44140 25596 44192
rect 25648 44180 25654 44192
rect 26421 44183 26479 44189
rect 26421 44180 26433 44183
rect 25648 44152 26433 44180
rect 25648 44140 25654 44152
rect 26421 44149 26433 44152
rect 26467 44149 26479 44183
rect 26421 44143 26479 44149
rect 27338 44140 27344 44192
rect 27396 44140 27402 44192
rect 28077 44183 28135 44189
rect 28077 44149 28089 44183
rect 28123 44180 28135 44183
rect 28718 44180 28724 44192
rect 28123 44152 28724 44180
rect 28123 44149 28135 44152
rect 28077 44143 28135 44149
rect 28718 44140 28724 44152
rect 28776 44140 28782 44192
rect 29104 44189 29132 44220
rect 29178 44208 29184 44260
rect 29236 44208 29242 44260
rect 30193 44251 30251 44257
rect 30193 44248 30205 44251
rect 29288 44220 30205 44248
rect 29089 44183 29147 44189
rect 29089 44149 29101 44183
rect 29135 44180 29147 44183
rect 29288 44180 29316 44220
rect 30193 44217 30205 44220
rect 30239 44248 30251 44251
rect 30834 44248 30840 44260
rect 30239 44220 30840 44248
rect 30239 44217 30251 44220
rect 30193 44211 30251 44217
rect 30834 44208 30840 44220
rect 30892 44208 30898 44260
rect 34793 44251 34851 44257
rect 34793 44217 34805 44251
rect 34839 44248 34851 44251
rect 35253 44251 35311 44257
rect 35253 44248 35265 44251
rect 34839 44220 35265 44248
rect 34839 44217 34851 44220
rect 34793 44211 34851 44217
rect 35253 44217 35265 44220
rect 35299 44217 35311 44251
rect 35253 44211 35311 44217
rect 37384 44220 37688 44248
rect 29135 44152 29316 44180
rect 29135 44149 29147 44152
rect 29089 44143 29147 44149
rect 29362 44140 29368 44192
rect 29420 44140 29426 44192
rect 30742 44140 30748 44192
rect 30800 44180 30806 44192
rect 31113 44183 31171 44189
rect 31113 44180 31125 44183
rect 30800 44152 31125 44180
rect 30800 44140 30806 44152
rect 31113 44149 31125 44152
rect 31159 44149 31171 44183
rect 31113 44143 31171 44149
rect 32398 44140 32404 44192
rect 32456 44180 32462 44192
rect 32953 44183 33011 44189
rect 32953 44180 32965 44183
rect 32456 44152 32965 44180
rect 32456 44140 32462 44152
rect 32953 44149 32965 44152
rect 32999 44149 33011 44183
rect 32953 44143 33011 44149
rect 33318 44140 33324 44192
rect 33376 44140 33382 44192
rect 33410 44140 33416 44192
rect 33468 44140 33474 44192
rect 33962 44140 33968 44192
rect 34020 44180 34026 44192
rect 34425 44183 34483 44189
rect 34425 44180 34437 44183
rect 34020 44152 34437 44180
rect 34020 44140 34026 44152
rect 34425 44149 34437 44152
rect 34471 44149 34483 44183
rect 34425 44143 34483 44149
rect 34885 44183 34943 44189
rect 34885 44149 34897 44183
rect 34931 44180 34943 44183
rect 35526 44180 35532 44192
rect 34931 44152 35532 44180
rect 34931 44149 34943 44152
rect 34885 44143 34943 44149
rect 35526 44140 35532 44152
rect 35584 44140 35590 44192
rect 36630 44140 36636 44192
rect 36688 44180 36694 44192
rect 37384 44180 37412 44220
rect 36688 44152 37412 44180
rect 36688 44140 36694 44152
rect 37458 44140 37464 44192
rect 37516 44140 37522 44192
rect 37660 44180 37688 44220
rect 37734 44208 37740 44260
rect 37792 44248 37798 44260
rect 37921 44251 37979 44257
rect 37921 44248 37933 44251
rect 37792 44220 37933 44248
rect 37792 44208 37798 44220
rect 37921 44217 37933 44220
rect 37967 44217 37979 44251
rect 37921 44211 37979 44217
rect 38102 44208 38108 44260
rect 38160 44248 38166 44260
rect 38746 44248 38752 44260
rect 38160 44220 38752 44248
rect 38160 44208 38166 44220
rect 38746 44208 38752 44220
rect 38804 44248 38810 44260
rect 39301 44251 39359 44257
rect 39301 44248 39313 44251
rect 38804 44220 39313 44248
rect 38804 44208 38810 44220
rect 39301 44217 39313 44220
rect 39347 44217 39359 44251
rect 39301 44211 39359 44217
rect 39945 44251 40003 44257
rect 39945 44217 39957 44251
rect 39991 44217 40003 44251
rect 39945 44211 40003 44217
rect 38838 44180 38844 44192
rect 37660 44152 38844 44180
rect 38838 44140 38844 44152
rect 38896 44140 38902 44192
rect 38933 44183 38991 44189
rect 38933 44149 38945 44183
rect 38979 44180 38991 44183
rect 39022 44180 39028 44192
rect 38979 44152 39028 44180
rect 38979 44149 38991 44152
rect 38933 44143 38991 44149
rect 39022 44140 39028 44152
rect 39080 44140 39086 44192
rect 39574 44140 39580 44192
rect 39632 44180 39638 44192
rect 39960 44180 39988 44211
rect 40494 44208 40500 44260
rect 40552 44248 40558 44260
rect 40681 44251 40739 44257
rect 40681 44248 40693 44251
rect 40552 44220 40693 44248
rect 40552 44208 40558 44220
rect 40681 44217 40693 44220
rect 40727 44217 40739 44251
rect 40681 44211 40739 44217
rect 40862 44208 40868 44260
rect 40920 44248 40926 44260
rect 41233 44251 41291 44257
rect 41233 44248 41245 44251
rect 40920 44220 41245 44248
rect 40920 44208 40926 44220
rect 41233 44217 41245 44220
rect 41279 44217 41291 44251
rect 41233 44211 41291 44217
rect 41340 44180 41368 44288
rect 43806 44276 43812 44328
rect 43864 44316 43870 44328
rect 44085 44319 44143 44325
rect 44085 44316 44097 44319
rect 43864 44288 44097 44316
rect 43864 44276 43870 44288
rect 44085 44285 44097 44288
rect 44131 44285 44143 44319
rect 46400 44316 46428 44424
rect 46753 44387 46811 44393
rect 46753 44353 46765 44387
rect 46799 44384 46811 44387
rect 48133 44387 48191 44393
rect 48133 44384 48145 44387
rect 46799 44356 48145 44384
rect 46799 44353 46811 44356
rect 46753 44347 46811 44353
rect 48133 44353 48145 44356
rect 48179 44384 48191 44387
rect 48222 44384 48228 44396
rect 48179 44356 48228 44384
rect 48179 44353 48191 44356
rect 48133 44347 48191 44353
rect 48222 44344 48228 44356
rect 48280 44344 48286 44396
rect 46400 44288 47348 44316
rect 44085 44279 44143 44285
rect 43073 44251 43131 44257
rect 43073 44217 43085 44251
rect 43119 44248 43131 44251
rect 43533 44251 43591 44257
rect 43533 44248 43545 44251
rect 43119 44220 43545 44248
rect 43119 44217 43131 44220
rect 43073 44211 43131 44217
rect 43533 44217 43545 44220
rect 43579 44217 43591 44251
rect 43533 44211 43591 44217
rect 46477 44251 46535 44257
rect 46477 44217 46489 44251
rect 46523 44248 46535 44251
rect 47029 44251 47087 44257
rect 47029 44248 47041 44251
rect 46523 44220 47041 44248
rect 46523 44217 46535 44220
rect 46477 44211 46535 44217
rect 47029 44217 47041 44220
rect 47075 44217 47087 44251
rect 47320 44248 47348 44288
rect 47394 44276 47400 44328
rect 47452 44316 47458 44328
rect 47581 44319 47639 44325
rect 47581 44316 47593 44319
rect 47452 44288 47593 44316
rect 47452 44276 47458 44288
rect 47581 44285 47593 44288
rect 47627 44285 47639 44319
rect 47581 44279 47639 44285
rect 47857 44251 47915 44257
rect 47857 44248 47869 44251
rect 47320 44220 47869 44248
rect 47029 44211 47087 44217
rect 47857 44217 47869 44220
rect 47903 44248 47915 44251
rect 50338 44248 50344 44260
rect 47903 44220 50344 44248
rect 47903 44217 47915 44220
rect 47857 44211 47915 44217
rect 50338 44208 50344 44220
rect 50396 44208 50402 44260
rect 39632 44152 41368 44180
rect 39632 44140 39638 44152
rect 41506 44140 41512 44192
rect 41564 44180 41570 44192
rect 41877 44183 41935 44189
rect 41877 44180 41889 44183
rect 41564 44152 41889 44180
rect 41564 44140 41570 44152
rect 41877 44149 41889 44152
rect 41923 44149 41935 44183
rect 41877 44143 41935 44149
rect 42242 44140 42248 44192
rect 42300 44140 42306 44192
rect 42334 44140 42340 44192
rect 42392 44140 42398 44192
rect 42426 44140 42432 44192
rect 42484 44180 42490 44192
rect 42705 44183 42763 44189
rect 42705 44180 42717 44183
rect 42484 44152 42717 44180
rect 42484 44140 42490 44152
rect 42705 44149 42717 44152
rect 42751 44149 42763 44183
rect 42705 44143 42763 44149
rect 43165 44183 43223 44189
rect 43165 44149 43177 44183
rect 43211 44180 43223 44183
rect 44450 44180 44456 44192
rect 43211 44152 44456 44180
rect 43211 44149 43223 44152
rect 43165 44143 43223 44149
rect 44450 44140 44456 44152
rect 44508 44140 44514 44192
rect 45370 44140 45376 44192
rect 45428 44180 45434 44192
rect 46109 44183 46167 44189
rect 46109 44180 46121 44183
rect 45428 44152 46121 44180
rect 45428 44140 45434 44152
rect 46109 44149 46121 44152
rect 46155 44149 46167 44183
rect 46109 44143 46167 44149
rect 46569 44183 46627 44189
rect 46569 44149 46581 44183
rect 46615 44180 46627 44183
rect 46934 44180 46940 44192
rect 46615 44152 46940 44180
rect 46615 44149 46627 44152
rect 46569 44143 46627 44149
rect 46934 44140 46940 44152
rect 46992 44140 46998 44192
rect 552 44090 66424 44112
rect 552 44038 2918 44090
rect 2970 44038 2982 44090
rect 3034 44038 3046 44090
rect 3098 44038 3110 44090
rect 3162 44038 3174 44090
rect 3226 44038 51918 44090
rect 51970 44038 51982 44090
rect 52034 44038 52046 44090
rect 52098 44038 52110 44090
rect 52162 44038 52174 44090
rect 52226 44038 66424 44090
rect 552 44016 66424 44038
rect 11606 43936 11612 43988
rect 11664 43976 11670 43988
rect 11977 43979 12035 43985
rect 11977 43976 11989 43979
rect 11664 43948 11989 43976
rect 11664 43936 11670 43948
rect 11977 43945 11989 43948
rect 12023 43945 12035 43979
rect 11977 43939 12035 43945
rect 14366 43936 14372 43988
rect 14424 43936 14430 43988
rect 14826 43936 14832 43988
rect 14884 43936 14890 43988
rect 16114 43936 16120 43988
rect 16172 43976 16178 43988
rect 19797 43979 19855 43985
rect 16172 43948 19380 43976
rect 16172 43936 16178 43948
rect 12986 43868 12992 43920
rect 13044 43908 13050 43920
rect 16485 43911 16543 43917
rect 13044 43880 13386 43908
rect 13044 43868 13050 43880
rect 16485 43877 16497 43911
rect 16531 43908 16543 43911
rect 16850 43908 16856 43920
rect 16531 43880 16856 43908
rect 16531 43877 16543 43880
rect 16485 43871 16543 43877
rect 16850 43868 16856 43880
rect 16908 43868 16914 43920
rect 17310 43868 17316 43920
rect 17368 43868 17374 43920
rect 17494 43868 17500 43920
rect 17552 43908 17558 43920
rect 17552 43880 17894 43908
rect 17552 43868 17558 43880
rect 18966 43868 18972 43920
rect 19024 43908 19030 43920
rect 19061 43911 19119 43917
rect 19061 43908 19073 43911
rect 19024 43880 19073 43908
rect 19024 43868 19030 43880
rect 19061 43877 19073 43880
rect 19107 43877 19119 43911
rect 19061 43871 19119 43877
rect 19352 43908 19380 43948
rect 19797 43945 19809 43979
rect 19843 43976 19855 43979
rect 20257 43979 20315 43985
rect 20257 43976 20269 43979
rect 19843 43948 20269 43976
rect 19843 43945 19855 43948
rect 19797 43939 19855 43945
rect 20257 43945 20269 43948
rect 20303 43945 20315 43979
rect 20257 43939 20315 43945
rect 24118 43936 24124 43988
rect 24176 43976 24182 43988
rect 24176 43948 25636 43976
rect 24176 43936 24182 43948
rect 20714 43908 20720 43920
rect 19352 43880 20720 43908
rect 11146 43800 11152 43852
rect 11204 43800 11210 43852
rect 12069 43843 12127 43849
rect 12069 43809 12081 43843
rect 12115 43840 12127 43843
rect 12526 43840 12532 43852
rect 12115 43812 12532 43840
rect 12115 43809 12127 43812
rect 12069 43803 12127 43809
rect 12526 43800 12532 43812
rect 12584 43800 12590 43852
rect 14734 43800 14740 43852
rect 14792 43840 14798 43852
rect 14792 43812 15056 43840
rect 14792 43800 14798 43812
rect 12253 43775 12311 43781
rect 12253 43741 12265 43775
rect 12299 43741 12311 43775
rect 12434 43772 12440 43784
rect 12253 43735 12311 43741
rect 12268 43704 12296 43735
rect 12406 43732 12440 43772
rect 12492 43732 12498 43784
rect 15028 43781 15056 43812
rect 15286 43800 15292 43852
rect 15344 43800 15350 43852
rect 15654 43800 15660 43852
rect 15712 43800 15718 43852
rect 19352 43849 19380 43880
rect 20714 43868 20720 43880
rect 20772 43868 20778 43920
rect 21542 43868 21548 43920
rect 21600 43868 21606 43920
rect 22186 43868 22192 43920
rect 22244 43868 22250 43920
rect 24946 43868 24952 43920
rect 25004 43868 25010 43920
rect 25608 43908 25636 43948
rect 26234 43936 26240 43988
rect 26292 43976 26298 43988
rect 26878 43976 26884 43988
rect 26292 43948 26884 43976
rect 26292 43936 26298 43948
rect 26878 43936 26884 43948
rect 26936 43976 26942 43988
rect 36630 43976 36636 43988
rect 26936 43948 29408 43976
rect 26936 43936 26942 43948
rect 25608 43880 27200 43908
rect 16577 43843 16635 43849
rect 16577 43809 16589 43843
rect 16623 43840 16635 43843
rect 19337 43843 19395 43849
rect 16623 43812 17632 43840
rect 16623 43809 16635 43812
rect 16577 43803 16635 43809
rect 12621 43775 12679 43781
rect 12621 43741 12633 43775
rect 12667 43772 12679 43775
rect 12897 43775 12955 43781
rect 12667 43744 12756 43772
rect 12667 43741 12679 43744
rect 12621 43735 12679 43741
rect 12406 43704 12434 43732
rect 12268 43676 12434 43704
rect 12728 43648 12756 43744
rect 12897 43741 12909 43775
rect 12943 43772 12955 43775
rect 14921 43775 14979 43781
rect 12943 43744 14504 43772
rect 12943 43741 12955 43744
rect 12897 43735 12955 43741
rect 14476 43713 14504 43744
rect 14921 43741 14933 43775
rect 14967 43741 14979 43775
rect 14921 43735 14979 43741
rect 15013 43775 15071 43781
rect 15013 43741 15025 43775
rect 15059 43741 15071 43775
rect 15013 43735 15071 43741
rect 14461 43707 14519 43713
rect 14461 43673 14473 43707
rect 14507 43673 14519 43707
rect 14936 43704 14964 43735
rect 16390 43732 16396 43784
rect 16448 43772 16454 43784
rect 16761 43775 16819 43781
rect 16761 43772 16773 43775
rect 16448 43744 16773 43772
rect 16448 43732 16454 43744
rect 16761 43741 16773 43744
rect 16807 43772 16819 43775
rect 17037 43775 17095 43781
rect 17037 43772 17049 43775
rect 16807 43744 17049 43772
rect 16807 43741 16819 43744
rect 16761 43735 16819 43741
rect 17037 43741 17049 43744
rect 17083 43741 17095 43775
rect 17604 43772 17632 43812
rect 19337 43809 19349 43843
rect 19383 43809 19395 43843
rect 19337 43803 19395 43809
rect 19518 43800 19524 43852
rect 19576 43840 19582 43852
rect 19576 43812 20760 43840
rect 19576 43800 19582 43812
rect 19794 43772 19800 43784
rect 17604 43744 19800 43772
rect 17037 43735 17095 43741
rect 19794 43732 19800 43744
rect 19852 43732 19858 43784
rect 19886 43732 19892 43784
rect 19944 43732 19950 43784
rect 20073 43775 20131 43781
rect 20073 43741 20085 43775
rect 20119 43772 20131 43775
rect 20622 43772 20628 43784
rect 20119 43744 20628 43772
rect 20119 43741 20131 43744
rect 20073 43735 20131 43741
rect 20622 43732 20628 43744
rect 20680 43732 20686 43784
rect 20732 43772 20760 43812
rect 20806 43800 20812 43852
rect 20864 43800 20870 43852
rect 22830 43800 22836 43852
rect 22888 43840 22894 43852
rect 23382 43840 23388 43852
rect 22888 43812 23388 43840
rect 22888 43800 22894 43812
rect 23382 43800 23388 43812
rect 23440 43840 23446 43852
rect 23477 43843 23535 43849
rect 23477 43840 23489 43843
rect 23440 43812 23489 43840
rect 23440 43800 23446 43812
rect 23477 43809 23489 43812
rect 23523 43809 23535 43843
rect 23477 43803 23535 43809
rect 26234 43800 26240 43852
rect 26292 43800 26298 43852
rect 27172 43849 27200 43880
rect 27338 43868 27344 43920
rect 27396 43868 27402 43920
rect 27706 43908 27712 43920
rect 27448 43880 27712 43908
rect 27157 43843 27215 43849
rect 27157 43809 27169 43843
rect 27203 43840 27215 43843
rect 27448 43840 27476 43880
rect 27706 43868 27712 43880
rect 27764 43868 27770 43920
rect 27203 43812 27476 43840
rect 27203 43809 27215 43812
rect 27157 43803 27215 43809
rect 28902 43800 28908 43852
rect 28960 43800 28966 43852
rect 29380 43849 29408 43948
rect 31726 43948 36636 43976
rect 29638 43868 29644 43920
rect 29696 43868 29702 43920
rect 29365 43843 29423 43849
rect 29365 43809 29377 43843
rect 29411 43809 29423 43843
rect 29365 43803 29423 43809
rect 30650 43800 30656 43852
rect 30708 43840 30714 43852
rect 30708 43812 30774 43840
rect 30708 43800 30714 43812
rect 21269 43775 21327 43781
rect 21269 43772 21281 43775
rect 20732 43744 21281 43772
rect 21269 43741 21281 43744
rect 21315 43741 21327 43775
rect 21269 43735 21327 43741
rect 22278 43732 22284 43784
rect 22336 43772 22342 43784
rect 22738 43772 22744 43784
rect 22336 43744 22744 43772
rect 22336 43732 22342 43744
rect 22738 43732 22744 43744
rect 22796 43772 22802 43784
rect 23017 43775 23075 43781
rect 23017 43772 23029 43775
rect 22796 43744 23029 43772
rect 22796 43732 22802 43744
rect 23017 43741 23029 43744
rect 23063 43741 23075 43775
rect 23017 43735 23075 43741
rect 23845 43775 23903 43781
rect 23845 43741 23857 43775
rect 23891 43772 23903 43775
rect 24489 43775 24547 43781
rect 24489 43772 24501 43775
rect 23891 43744 24501 43772
rect 23891 43741 23903 43744
rect 23845 43735 23903 43741
rect 24489 43741 24501 43744
rect 24535 43772 24547 43775
rect 25314 43772 25320 43784
rect 24535 43744 25320 43772
rect 24535 43741 24547 43744
rect 24489 43735 24547 43741
rect 25314 43732 25320 43744
rect 25372 43732 25378 43784
rect 25958 43732 25964 43784
rect 26016 43732 26022 43784
rect 26326 43732 26332 43784
rect 26384 43772 26390 43784
rect 26973 43775 27031 43781
rect 26973 43772 26985 43775
rect 26384 43744 26985 43772
rect 26384 43732 26390 43744
rect 26973 43741 26985 43744
rect 27019 43741 27031 43775
rect 26973 43735 27031 43741
rect 27062 43732 27068 43784
rect 27120 43772 27126 43784
rect 27525 43775 27583 43781
rect 27525 43772 27537 43775
rect 27120 43744 27537 43772
rect 27120 43732 27126 43744
rect 27525 43741 27537 43744
rect 27571 43741 27583 43775
rect 27525 43735 27583 43741
rect 27801 43775 27859 43781
rect 27801 43741 27813 43775
rect 27847 43772 27859 43775
rect 28994 43772 29000 43784
rect 27847 43744 29000 43772
rect 27847 43741 27859 43744
rect 27801 43735 27859 43741
rect 28994 43732 29000 43744
rect 29052 43732 29058 43784
rect 29273 43775 29331 43781
rect 29273 43741 29285 43775
rect 29319 43772 29331 43775
rect 30374 43772 30380 43784
rect 29319 43744 30380 43772
rect 29319 43741 29331 43744
rect 29273 43735 29331 43741
rect 30374 43732 30380 43744
rect 30432 43732 30438 43784
rect 31386 43732 31392 43784
rect 31444 43732 31450 43784
rect 16117 43707 16175 43713
rect 16117 43704 16129 43707
rect 14936 43676 16129 43704
rect 14461 43667 14519 43673
rect 16117 43673 16129 43676
rect 16163 43673 16175 43707
rect 17954 43704 17960 43716
rect 16117 43667 16175 43673
rect 16960 43676 17960 43704
rect 11054 43596 11060 43648
rect 11112 43636 11118 43648
rect 11609 43639 11667 43645
rect 11609 43636 11621 43639
rect 11112 43608 11621 43636
rect 11112 43596 11118 43608
rect 11609 43605 11621 43608
rect 11655 43605 11667 43639
rect 11609 43599 11667 43605
rect 12710 43596 12716 43648
rect 12768 43636 12774 43648
rect 14734 43636 14740 43648
rect 12768 43608 14740 43636
rect 12768 43596 12774 43608
rect 14734 43596 14740 43608
rect 14792 43596 14798 43648
rect 15841 43639 15899 43645
rect 15841 43605 15853 43639
rect 15887 43636 15899 43639
rect 16960 43636 16988 43676
rect 17954 43664 17960 43676
rect 18012 43664 18018 43716
rect 24397 43707 24455 43713
rect 24397 43673 24409 43707
rect 24443 43704 24455 43707
rect 24578 43704 24584 43716
rect 24443 43676 24584 43704
rect 24443 43673 24455 43676
rect 24397 43667 24455 43673
rect 24578 43664 24584 43676
rect 24636 43664 24642 43716
rect 31726 43704 31754 43948
rect 36630 43936 36636 43948
rect 36688 43936 36694 43988
rect 36725 43979 36783 43985
rect 36725 43945 36737 43979
rect 36771 43976 36783 43979
rect 37274 43976 37280 43988
rect 36771 43948 37280 43976
rect 36771 43945 36783 43948
rect 36725 43939 36783 43945
rect 37274 43936 37280 43948
rect 37332 43976 37338 43988
rect 38286 43976 38292 43988
rect 37332 43948 38292 43976
rect 37332 43936 37338 43948
rect 38286 43936 38292 43948
rect 38344 43936 38350 43988
rect 38838 43936 38844 43988
rect 38896 43976 38902 43988
rect 39761 43979 39819 43985
rect 39761 43976 39773 43979
rect 38896 43948 39773 43976
rect 38896 43936 38902 43948
rect 39761 43945 39773 43948
rect 39807 43976 39819 43979
rect 41046 43976 41052 43988
rect 39807 43948 41052 43976
rect 39807 43945 39819 43948
rect 39761 43939 39819 43945
rect 41046 43936 41052 43948
rect 41104 43936 41110 43988
rect 42242 43936 42248 43988
rect 42300 43976 42306 43988
rect 43901 43979 43959 43985
rect 43901 43976 43913 43979
rect 42300 43948 43913 43976
rect 42300 43936 42306 43948
rect 43901 43945 43913 43948
rect 43947 43945 43959 43979
rect 43901 43939 43959 43945
rect 46845 43979 46903 43985
rect 46845 43945 46857 43979
rect 46891 43976 46903 43979
rect 47394 43976 47400 43988
rect 46891 43948 47400 43976
rect 46891 43945 46903 43948
rect 46845 43939 46903 43945
rect 47394 43936 47400 43948
rect 47452 43936 47458 43988
rect 33962 43868 33968 43920
rect 34020 43868 34026 43920
rect 34054 43868 34060 43920
rect 34112 43908 34118 43920
rect 38102 43908 38108 43920
rect 34112 43880 34454 43908
rect 37766 43880 38108 43908
rect 34112 43868 34118 43880
rect 38102 43868 38108 43880
rect 38160 43868 38166 43920
rect 38197 43911 38255 43917
rect 38197 43877 38209 43911
rect 38243 43908 38255 43911
rect 38654 43908 38660 43920
rect 38243 43880 38660 43908
rect 38243 43877 38255 43880
rect 38197 43871 38255 43877
rect 38654 43868 38660 43880
rect 38712 43868 38718 43920
rect 42337 43911 42395 43917
rect 38856 43880 39896 43908
rect 31846 43800 31852 43852
rect 31904 43800 31910 43852
rect 32769 43843 32827 43849
rect 32769 43809 32781 43843
rect 32815 43840 32827 43843
rect 33229 43843 33287 43849
rect 33229 43840 33241 43843
rect 32815 43812 33241 43840
rect 32815 43809 32827 43812
rect 32769 43803 32827 43809
rect 33229 43809 33241 43812
rect 33275 43809 33287 43843
rect 33229 43803 33287 43809
rect 35897 43843 35955 43849
rect 35897 43809 35909 43843
rect 35943 43840 35955 43843
rect 36630 43840 36636 43852
rect 35943 43812 36636 43840
rect 35943 43809 35955 43812
rect 35897 43803 35955 43809
rect 36630 43800 36636 43812
rect 36688 43800 36694 43852
rect 38473 43843 38531 43849
rect 38473 43809 38485 43843
rect 38519 43840 38531 43843
rect 38856 43840 38884 43880
rect 38519 43812 38884 43840
rect 38519 43809 38531 43812
rect 38473 43803 38531 43809
rect 38930 43800 38936 43852
rect 38988 43800 38994 43852
rect 39390 43800 39396 43852
rect 39448 43800 39454 43852
rect 32214 43732 32220 43784
rect 32272 43732 32278 43784
rect 33042 43732 33048 43784
rect 33100 43732 33106 43784
rect 33137 43775 33195 43781
rect 33137 43741 33149 43775
rect 33183 43772 33195 43775
rect 33594 43772 33600 43784
rect 33183 43744 33600 43772
rect 33183 43741 33195 43744
rect 33137 43735 33195 43741
rect 33594 43732 33600 43744
rect 33652 43732 33658 43784
rect 33689 43775 33747 43781
rect 33689 43741 33701 43775
rect 33735 43741 33747 43775
rect 33689 43735 33747 43741
rect 30668 43676 31754 43704
rect 15887 43608 16988 43636
rect 17589 43639 17647 43645
rect 15887 43605 15899 43608
rect 15841 43599 15899 43605
rect 17589 43605 17601 43639
rect 17635 43636 17647 43639
rect 18046 43636 18052 43648
rect 17635 43608 18052 43636
rect 17635 43605 17647 43608
rect 17589 43599 17647 43605
rect 18046 43596 18052 43608
rect 18104 43636 18110 43648
rect 19242 43636 19248 43648
rect 18104 43608 19248 43636
rect 18104 43596 18110 43608
rect 19242 43596 19248 43608
rect 19300 43596 19306 43648
rect 19426 43596 19432 43648
rect 19484 43596 19490 43648
rect 20070 43596 20076 43648
rect 20128 43636 20134 43648
rect 21910 43636 21916 43648
rect 20128 43608 21916 43636
rect 20128 43596 20134 43608
rect 21910 43596 21916 43608
rect 21968 43596 21974 43648
rect 22646 43596 22652 43648
rect 22704 43636 22710 43648
rect 23201 43639 23259 43645
rect 23201 43636 23213 43639
rect 22704 43608 23213 43636
rect 22704 43596 22710 43608
rect 23201 43605 23213 43608
rect 23247 43605 23259 43639
rect 23201 43599 23259 43605
rect 26234 43596 26240 43648
rect 26292 43636 26298 43648
rect 26421 43639 26479 43645
rect 26421 43636 26433 43639
rect 26292 43608 26433 43636
rect 26292 43596 26298 43608
rect 26421 43605 26433 43608
rect 26467 43605 26479 43639
rect 26421 43599 26479 43605
rect 26510 43596 26516 43648
rect 26568 43636 26574 43648
rect 30668 43636 30696 43676
rect 32122 43664 32128 43716
rect 32180 43704 32186 43716
rect 33704 43704 33732 43735
rect 35434 43732 35440 43784
rect 35492 43732 35498 43784
rect 35989 43775 36047 43781
rect 35989 43772 36001 43775
rect 35866 43744 36001 43772
rect 32180 43676 33732 43704
rect 32180 43664 32186 43676
rect 35526 43664 35532 43716
rect 35584 43664 35590 43716
rect 26568 43608 30696 43636
rect 26568 43596 26574 43608
rect 31662 43596 31668 43648
rect 31720 43636 31726 43648
rect 33226 43636 33232 43648
rect 31720 43608 33232 43636
rect 31720 43596 31726 43608
rect 33226 43596 33232 43608
rect 33284 43596 33290 43648
rect 33597 43639 33655 43645
rect 33597 43605 33609 43639
rect 33643 43636 33655 43639
rect 33686 43636 33692 43648
rect 33643 43608 33692 43636
rect 33643 43605 33655 43608
rect 33597 43599 33655 43605
rect 33686 43596 33692 43608
rect 33744 43596 33750 43648
rect 34330 43596 34336 43648
rect 34388 43636 34394 43648
rect 35866 43636 35894 43744
rect 35989 43741 36001 43744
rect 36035 43741 36047 43775
rect 35989 43735 36047 43741
rect 36173 43775 36231 43781
rect 36173 43741 36185 43775
rect 36219 43772 36231 43775
rect 37550 43772 37556 43784
rect 36219 43744 37556 43772
rect 36219 43741 36231 43744
rect 36173 43735 36231 43741
rect 37550 43732 37556 43744
rect 37608 43772 37614 43784
rect 38657 43775 38715 43781
rect 38657 43772 38669 43775
rect 37608 43744 38669 43772
rect 37608 43732 37614 43744
rect 38657 43741 38669 43744
rect 38703 43741 38715 43775
rect 38657 43735 38715 43741
rect 38841 43775 38899 43781
rect 38841 43741 38853 43775
rect 38887 43741 38899 43775
rect 39868 43772 39896 43880
rect 42337 43877 42349 43911
rect 42383 43908 42395 43911
rect 42426 43908 42432 43920
rect 42383 43880 42432 43908
rect 42383 43877 42395 43880
rect 42337 43871 42395 43877
rect 42426 43868 42432 43880
rect 42484 43868 42490 43920
rect 42886 43868 42892 43920
rect 42944 43868 42950 43920
rect 45370 43868 45376 43920
rect 45428 43868 45434 43920
rect 46014 43868 46020 43920
rect 46072 43868 46078 43920
rect 39942 43800 39948 43852
rect 40000 43840 40006 43852
rect 44453 43843 44511 43849
rect 44453 43840 44465 43843
rect 40000 43812 40158 43840
rect 43548 43812 44465 43840
rect 40000 43800 40006 43812
rect 40218 43772 40224 43784
rect 39868 43744 40224 43772
rect 38841 43735 38899 43741
rect 34388 43608 35894 43636
rect 34388 43596 34394 43608
rect 36630 43596 36636 43648
rect 36688 43636 36694 43648
rect 38856 43636 38884 43735
rect 40218 43732 40224 43744
rect 40276 43772 40282 43784
rect 40770 43772 40776 43784
rect 40276 43744 40776 43772
rect 40276 43732 40282 43744
rect 40770 43732 40776 43744
rect 40828 43732 40834 43784
rect 41233 43775 41291 43781
rect 41233 43741 41245 43775
rect 41279 43772 41291 43775
rect 41509 43775 41567 43781
rect 41279 43744 41460 43772
rect 41279 43741 41291 43744
rect 41233 43735 41291 43741
rect 39574 43664 39580 43716
rect 39632 43664 39638 43716
rect 41432 43648 41460 43744
rect 41509 43741 41521 43775
rect 41555 43772 41567 43775
rect 41966 43772 41972 43784
rect 41555 43744 41972 43772
rect 41555 43741 41567 43744
rect 41509 43735 41567 43741
rect 41966 43732 41972 43744
rect 42024 43772 42030 43784
rect 42061 43775 42119 43781
rect 42061 43772 42073 43775
rect 42024 43744 42073 43772
rect 42024 43732 42030 43744
rect 42061 43741 42073 43744
rect 42107 43741 42119 43775
rect 42061 43735 42119 43741
rect 42702 43732 42708 43784
rect 42760 43772 42766 43784
rect 43548 43772 43576 43812
rect 44453 43809 44465 43812
rect 44499 43809 44511 43843
rect 44453 43803 44511 43809
rect 48038 43800 48044 43852
rect 48096 43840 48102 43852
rect 48225 43843 48283 43849
rect 48225 43840 48237 43843
rect 48096 43812 48237 43840
rect 48096 43800 48102 43812
rect 48225 43809 48237 43812
rect 48271 43809 48283 43843
rect 48225 43803 48283 43809
rect 42760 43744 43576 43772
rect 42760 43732 42766 43744
rect 43806 43732 43812 43784
rect 43864 43732 43870 43784
rect 45094 43732 45100 43784
rect 45152 43732 45158 43784
rect 47210 43732 47216 43784
rect 47268 43772 47274 43784
rect 47489 43775 47547 43781
rect 47489 43772 47501 43775
rect 47268 43744 47501 43772
rect 47268 43732 47274 43744
rect 47489 43741 47501 43744
rect 47535 43741 47547 43775
rect 47489 43735 47547 43741
rect 47578 43732 47584 43784
rect 47636 43732 47642 43784
rect 48682 43732 48688 43784
rect 48740 43732 48746 43784
rect 36688 43608 38884 43636
rect 36688 43596 36694 43608
rect 39298 43596 39304 43648
rect 39356 43596 39362 43648
rect 41414 43596 41420 43648
rect 41472 43596 41478 43648
rect 47029 43639 47087 43645
rect 47029 43605 47041 43639
rect 47075 43636 47087 43639
rect 47302 43636 47308 43648
rect 47075 43608 47308 43636
rect 47075 43605 47087 43608
rect 47029 43599 47087 43605
rect 47302 43596 47308 43608
rect 47360 43596 47366 43648
rect 47762 43596 47768 43648
rect 47820 43636 47826 43648
rect 47949 43639 48007 43645
rect 47949 43636 47961 43639
rect 47820 43608 47961 43636
rect 47820 43596 47826 43608
rect 47949 43605 47961 43608
rect 47995 43605 48007 43639
rect 47949 43599 48007 43605
rect 49237 43639 49295 43645
rect 49237 43605 49249 43639
rect 49283 43636 49295 43639
rect 49418 43636 49424 43648
rect 49283 43608 49424 43636
rect 49283 43605 49295 43608
rect 49237 43599 49295 43605
rect 49418 43596 49424 43608
rect 49476 43596 49482 43648
rect 552 43546 66424 43568
rect 552 43494 1998 43546
rect 2050 43494 2062 43546
rect 2114 43494 2126 43546
rect 2178 43494 2190 43546
rect 2242 43494 2254 43546
rect 2306 43494 50998 43546
rect 51050 43494 51062 43546
rect 51114 43494 51126 43546
rect 51178 43494 51190 43546
rect 51242 43494 51254 43546
rect 51306 43494 66424 43546
rect 552 43472 66424 43494
rect 12710 43432 12716 43444
rect 11348 43404 12716 43432
rect 11054 43256 11060 43308
rect 11112 43256 11118 43308
rect 11348 43305 11376 43404
rect 12710 43392 12716 43404
rect 12768 43392 12774 43444
rect 13998 43392 14004 43444
rect 14056 43432 14062 43444
rect 15289 43435 15347 43441
rect 15289 43432 15301 43435
rect 14056 43404 15301 43432
rect 14056 43392 14062 43404
rect 15289 43401 15301 43404
rect 15335 43432 15347 43435
rect 16850 43432 16856 43444
rect 15335 43404 16856 43432
rect 15335 43401 15347 43404
rect 15289 43395 15347 43401
rect 16850 43392 16856 43404
rect 16908 43392 16914 43444
rect 16942 43392 16948 43444
rect 17000 43432 17006 43444
rect 17494 43432 17500 43444
rect 17000 43404 17500 43432
rect 17000 43392 17006 43404
rect 17494 43392 17500 43404
rect 17552 43432 17558 43444
rect 19610 43432 19616 43444
rect 17552 43404 19616 43432
rect 17552 43392 17558 43404
rect 19610 43392 19616 43404
rect 19668 43392 19674 43444
rect 19797 43435 19855 43441
rect 19797 43401 19809 43435
rect 19843 43432 19855 43435
rect 19886 43432 19892 43444
rect 19843 43404 19892 43432
rect 19843 43401 19855 43404
rect 19797 43395 19855 43401
rect 19886 43392 19892 43404
rect 19944 43392 19950 43444
rect 20364 43404 21588 43432
rect 18782 43324 18788 43376
rect 18840 43324 18846 43376
rect 20364 43364 20392 43404
rect 19076 43336 20392 43364
rect 21560 43364 21588 43404
rect 21910 43392 21916 43444
rect 21968 43392 21974 43444
rect 22094 43392 22100 43444
rect 22152 43392 22158 43444
rect 23934 43392 23940 43444
rect 23992 43392 23998 43444
rect 25590 43432 25596 43444
rect 24044 43404 25596 43432
rect 23566 43364 23572 43376
rect 21560 43336 23572 43364
rect 19076 43308 19104 43336
rect 23566 43324 23572 43336
rect 23624 43324 23630 43376
rect 24044 43364 24072 43404
rect 25590 43392 25596 43404
rect 25648 43392 25654 43444
rect 25958 43392 25964 43444
rect 26016 43432 26022 43444
rect 26053 43435 26111 43441
rect 26053 43432 26065 43435
rect 26016 43404 26065 43432
rect 26016 43392 26022 43404
rect 26053 43401 26065 43404
rect 26099 43401 26111 43435
rect 26053 43395 26111 43401
rect 28626 43392 28632 43444
rect 28684 43392 28690 43444
rect 28994 43392 29000 43444
rect 29052 43392 29058 43444
rect 29638 43392 29644 43444
rect 29696 43432 29702 43444
rect 29825 43435 29883 43441
rect 29825 43432 29837 43435
rect 29696 43404 29837 43432
rect 29696 43392 29702 43404
rect 29825 43401 29837 43404
rect 29871 43401 29883 43435
rect 29825 43395 29883 43401
rect 30098 43392 30104 43444
rect 30156 43432 30162 43444
rect 31570 43432 31576 43444
rect 30156 43404 31576 43432
rect 30156 43392 30162 43404
rect 31570 43392 31576 43404
rect 31628 43432 31634 43444
rect 33134 43432 33140 43444
rect 31628 43404 33140 43432
rect 31628 43392 31634 43404
rect 33134 43392 33140 43404
rect 33192 43392 33198 43444
rect 33318 43392 33324 43444
rect 33376 43432 33382 43444
rect 34149 43435 34207 43441
rect 34149 43432 34161 43435
rect 33376 43404 34161 43432
rect 33376 43392 33382 43404
rect 34149 43401 34161 43404
rect 34195 43401 34207 43435
rect 34149 43395 34207 43401
rect 34238 43392 34244 43444
rect 34296 43432 34302 43444
rect 36538 43432 36544 43444
rect 34296 43404 36544 43432
rect 34296 43392 34302 43404
rect 36538 43392 36544 43404
rect 36596 43392 36602 43444
rect 36630 43392 36636 43444
rect 36688 43392 36694 43444
rect 37918 43392 37924 43444
rect 37976 43432 37982 43444
rect 39301 43435 39359 43441
rect 39301 43432 39313 43435
rect 37976 43404 39313 43432
rect 37976 43392 37982 43404
rect 39301 43401 39313 43404
rect 39347 43401 39359 43435
rect 39301 43395 39359 43401
rect 40126 43392 40132 43444
rect 40184 43432 40190 43444
rect 40313 43435 40371 43441
rect 40313 43432 40325 43435
rect 40184 43404 40325 43432
rect 40184 43392 40190 43404
rect 40313 43401 40325 43404
rect 40359 43432 40371 43435
rect 40359 43404 42288 43432
rect 40359 43401 40371 43404
rect 40313 43395 40371 43401
rect 23860 43336 24072 43364
rect 11333 43299 11391 43305
rect 11333 43265 11345 43299
rect 11379 43265 11391 43299
rect 11333 43259 11391 43265
rect 11425 43299 11483 43305
rect 11425 43265 11437 43299
rect 11471 43296 11483 43299
rect 13541 43299 13599 43305
rect 13541 43296 13553 43299
rect 11471 43268 13553 43296
rect 11471 43265 11483 43268
rect 11425 43259 11483 43265
rect 13541 43265 13553 43268
rect 13587 43296 13599 43299
rect 16114 43296 16120 43308
rect 13587 43268 16120 43296
rect 13587 43265 13599 43268
rect 13541 43259 13599 43265
rect 16114 43256 16120 43268
rect 16172 43256 16178 43308
rect 19058 43256 19064 43308
rect 19116 43256 19122 43308
rect 19153 43299 19211 43305
rect 19153 43265 19165 43299
rect 19199 43296 19211 43299
rect 19334 43296 19340 43308
rect 19199 43268 19340 43296
rect 19199 43265 19211 43268
rect 19153 43259 19211 43265
rect 19334 43256 19340 43268
rect 19392 43256 19398 43308
rect 19610 43256 19616 43308
rect 19668 43296 19674 43308
rect 20162 43296 20168 43308
rect 19668 43268 20168 43296
rect 19668 43256 19674 43268
rect 20162 43256 20168 43268
rect 20220 43256 20226 43308
rect 20714 43256 20720 43308
rect 20772 43296 20778 43308
rect 21637 43299 21695 43305
rect 21637 43296 21649 43299
rect 20772 43268 21649 43296
rect 20772 43256 20778 43268
rect 21637 43265 21649 43268
rect 21683 43265 21695 43299
rect 22462 43296 22468 43308
rect 21637 43259 21695 43265
rect 21836 43268 22468 43296
rect 16022 43188 16028 43240
rect 16080 43188 16086 43240
rect 16206 43188 16212 43240
rect 16264 43188 16270 43240
rect 18969 43231 19027 43237
rect 18969 43197 18981 43231
rect 19015 43197 19027 43231
rect 18969 43191 19027 43197
rect 10594 43120 10600 43172
rect 10652 43120 10658 43172
rect 11698 43120 11704 43172
rect 11756 43120 11762 43172
rect 12986 43160 12992 43172
rect 12926 43132 12992 43160
rect 12986 43120 12992 43132
rect 13044 43160 13050 43172
rect 13044 43132 13768 43160
rect 13044 43120 13050 43132
rect 9585 43095 9643 43101
rect 9585 43061 9597 43095
rect 9631 43092 9643 43095
rect 12342 43092 12348 43104
rect 9631 43064 12348 43092
rect 9631 43061 9643 43064
rect 9585 43055 9643 43061
rect 12342 43052 12348 43064
rect 12400 43052 12406 43104
rect 13170 43052 13176 43104
rect 13228 43052 13234 43104
rect 13740 43092 13768 43132
rect 13814 43120 13820 43172
rect 13872 43120 13878 43172
rect 14274 43160 14280 43172
rect 13924 43132 14280 43160
rect 13924 43092 13952 43132
rect 14274 43120 14280 43132
rect 14332 43120 14338 43172
rect 16485 43163 16543 43169
rect 16485 43129 16497 43163
rect 16531 43160 16543 43163
rect 16574 43160 16580 43172
rect 16531 43132 16580 43160
rect 16531 43129 16543 43132
rect 16485 43123 16543 43129
rect 16574 43120 16580 43132
rect 16632 43120 16638 43172
rect 16942 43120 16948 43172
rect 17000 43120 17006 43172
rect 18984 43160 19012 43191
rect 19242 43188 19248 43240
rect 19300 43228 19306 43240
rect 19429 43231 19487 43237
rect 19429 43228 19441 43231
rect 19300 43200 19441 43228
rect 19300 43188 19306 43200
rect 19429 43197 19441 43200
rect 19475 43197 19487 43231
rect 19429 43191 19487 43197
rect 21726 43188 21732 43240
rect 21784 43188 21790 43240
rect 19337 43163 19395 43169
rect 19337 43160 19349 43163
rect 18984 43132 19349 43160
rect 19337 43129 19349 43132
rect 19383 43160 19395 43163
rect 19383 43132 19932 43160
rect 19383 43129 19395 43132
rect 19337 43123 19395 43129
rect 13740 43064 13952 43092
rect 15473 43095 15531 43101
rect 15473 43061 15485 43095
rect 15519 43092 15531 43095
rect 15562 43092 15568 43104
rect 15519 43064 15568 43092
rect 15519 43061 15531 43064
rect 15473 43055 15531 43061
rect 15562 43052 15568 43064
rect 15620 43052 15626 43104
rect 17957 43095 18015 43101
rect 17957 43061 17969 43095
rect 18003 43092 18015 43095
rect 18506 43092 18512 43104
rect 18003 43064 18512 43092
rect 18003 43061 18015 43064
rect 17957 43055 18015 43061
rect 18506 43052 18512 43064
rect 18564 43092 18570 43104
rect 19150 43092 19156 43104
rect 18564 43064 19156 43092
rect 18564 43052 18570 43064
rect 19150 43052 19156 43064
rect 19208 43052 19214 43104
rect 19904 43101 19932 43132
rect 20070 43120 20076 43172
rect 20128 43160 20134 43172
rect 21361 43163 21419 43169
rect 20128 43132 20194 43160
rect 20128 43120 20134 43132
rect 21361 43129 21373 43163
rect 21407 43160 21419 43163
rect 21836 43160 21864 43268
rect 22462 43256 22468 43268
rect 22520 43256 22526 43308
rect 22646 43256 22652 43308
rect 22704 43256 22710 43308
rect 23860 43296 23888 43336
rect 25498 43324 25504 43376
rect 25556 43364 25562 43376
rect 26234 43364 26240 43376
rect 25556 43336 26240 43364
rect 25556 43324 25562 43336
rect 26234 43324 26240 43336
rect 26292 43324 26298 43376
rect 26326 43324 26332 43376
rect 26384 43364 26390 43376
rect 26384 43336 27752 43364
rect 26384 43324 26390 43336
rect 23492 43268 23888 43296
rect 22557 43231 22615 43237
rect 22557 43197 22569 43231
rect 22603 43228 22615 43231
rect 23492 43228 23520 43268
rect 24578 43256 24584 43308
rect 24636 43296 24642 43308
rect 26620 43305 26648 43336
rect 26605 43299 26663 43305
rect 24636 43268 26464 43296
rect 24636 43256 24642 43268
rect 22603 43200 23520 43228
rect 23569 43231 23627 43237
rect 22603 43197 22615 43200
rect 22557 43191 22615 43197
rect 23569 43197 23581 43231
rect 23615 43197 23627 43231
rect 23569 43191 23627 43197
rect 22094 43160 22100 43172
rect 21407 43132 21864 43160
rect 21928 43132 22100 43160
rect 21407 43129 21419 43132
rect 21361 43123 21419 43129
rect 19889 43095 19947 43101
rect 19889 43061 19901 43095
rect 19935 43092 19947 43095
rect 21928 43092 21956 43132
rect 22094 43120 22100 43132
rect 22152 43160 22158 43172
rect 22465 43163 22523 43169
rect 22465 43160 22477 43163
rect 22152 43132 22477 43160
rect 22152 43120 22158 43132
rect 22465 43129 22477 43132
rect 22511 43129 22523 43163
rect 22465 43123 22523 43129
rect 19935 43064 21956 43092
rect 19935 43061 19947 43064
rect 19889 43055 19947 43061
rect 22002 43052 22008 43104
rect 22060 43092 22066 43104
rect 22186 43092 22192 43104
rect 22060 43064 22192 43092
rect 22060 43052 22066 43064
rect 22186 43052 22192 43064
rect 22244 43052 22250 43104
rect 22922 43052 22928 43104
rect 22980 43052 22986 43104
rect 23584 43092 23612 43191
rect 23658 43188 23664 43240
rect 23716 43228 23722 43240
rect 24118 43228 24124 43240
rect 23716 43200 24124 43228
rect 23716 43188 23722 43200
rect 24118 43188 24124 43200
rect 24176 43188 24182 43240
rect 26436 43237 26464 43268
rect 26605 43265 26617 43299
rect 26651 43265 26663 43299
rect 27525 43299 27583 43305
rect 27525 43296 27537 43299
rect 26605 43259 26663 43265
rect 26712 43268 27537 43296
rect 24213 43231 24271 43237
rect 24213 43197 24225 43231
rect 24259 43197 24271 43231
rect 24213 43191 24271 43197
rect 26421 43231 26479 43237
rect 26421 43197 26433 43231
rect 26467 43197 26479 43231
rect 26421 43191 26479 43197
rect 23842 43120 23848 43172
rect 23900 43160 23906 43172
rect 24228 43160 24256 43191
rect 23900 43132 24256 43160
rect 24489 43163 24547 43169
rect 23900 43120 23906 43132
rect 24489 43129 24501 43163
rect 24535 43160 24547 43163
rect 24578 43160 24584 43172
rect 24535 43132 24584 43160
rect 24535 43129 24547 43132
rect 24489 43123 24547 43129
rect 24578 43120 24584 43132
rect 24636 43120 24642 43172
rect 24946 43120 24952 43172
rect 25004 43120 25010 43172
rect 26712 43160 26740 43268
rect 27525 43265 27537 43268
rect 27571 43265 27583 43299
rect 27525 43259 27583 43265
rect 27614 43256 27620 43308
rect 27672 43256 27678 43308
rect 27724 43296 27752 43336
rect 28258 43324 28264 43376
rect 28316 43364 28322 43376
rect 28902 43364 28908 43376
rect 28316 43336 28908 43364
rect 28316 43324 28322 43336
rect 28902 43324 28908 43336
rect 28960 43364 28966 43376
rect 30742 43364 30748 43376
rect 28960 43336 30748 43364
rect 28960 43324 28966 43336
rect 30742 43324 30748 43336
rect 30800 43324 30806 43376
rect 28350 43296 28356 43308
rect 27724 43268 28356 43296
rect 28350 43256 28356 43268
rect 28408 43296 28414 43308
rect 29638 43296 29644 43308
rect 28408 43268 29644 43296
rect 28408 43256 28414 43268
rect 29638 43256 29644 43268
rect 29696 43256 29702 43308
rect 30098 43256 30104 43308
rect 30156 43296 30162 43308
rect 30377 43299 30435 43305
rect 30377 43296 30389 43299
rect 30156 43268 30389 43296
rect 30156 43256 30162 43268
rect 30377 43265 30389 43268
rect 30423 43265 30435 43299
rect 30377 43259 30435 43265
rect 33686 43256 33692 43308
rect 33744 43256 33750 43308
rect 33965 43299 34023 43305
rect 33965 43265 33977 43299
rect 34011 43296 34023 43299
rect 34885 43299 34943 43305
rect 34885 43296 34897 43299
rect 34011 43268 34897 43296
rect 34011 43265 34023 43268
rect 33965 43259 34023 43265
rect 34885 43265 34897 43268
rect 34931 43296 34943 43299
rect 37090 43296 37096 43308
rect 34931 43268 37096 43296
rect 34931 43265 34943 43268
rect 34885 43259 34943 43265
rect 37090 43256 37096 43268
rect 37148 43296 37154 43308
rect 37185 43299 37243 43305
rect 37185 43296 37197 43299
rect 37148 43268 37197 43296
rect 37148 43256 37154 43268
rect 37185 43265 37197 43268
rect 37231 43265 37243 43299
rect 37185 43259 37243 43265
rect 37458 43256 37464 43308
rect 37516 43256 37522 43308
rect 38930 43256 38936 43308
rect 38988 43256 38994 43308
rect 40770 43256 40776 43308
rect 40828 43296 40834 43308
rect 40957 43299 41015 43305
rect 40957 43296 40969 43299
rect 40828 43268 40969 43296
rect 40828 43256 40834 43268
rect 40957 43265 40969 43268
rect 41003 43296 41015 43299
rect 41322 43296 41328 43308
rect 41003 43268 41328 43296
rect 41003 43265 41015 43268
rect 40957 43259 41015 43265
rect 41322 43256 41328 43268
rect 41380 43256 41386 43308
rect 42260 43296 42288 43404
rect 42334 43392 42340 43444
rect 42392 43432 42398 43444
rect 42797 43435 42855 43441
rect 42797 43432 42809 43435
rect 42392 43404 42809 43432
rect 42392 43392 42398 43404
rect 42797 43401 42809 43404
rect 42843 43401 42855 43435
rect 42797 43395 42855 43401
rect 43070 43392 43076 43444
rect 43128 43432 43134 43444
rect 43128 43404 45048 43432
rect 43128 43392 43134 43404
rect 42702 43324 42708 43376
rect 42760 43324 42766 43376
rect 43806 43364 43812 43376
rect 43272 43336 43812 43364
rect 42610 43296 42616 43308
rect 42260 43268 42616 43296
rect 42610 43256 42616 43268
rect 42668 43296 42674 43308
rect 43272 43305 43300 43336
rect 43806 43324 43812 43336
rect 43864 43324 43870 43376
rect 45020 43305 45048 43404
rect 43257 43299 43315 43305
rect 42668 43268 43208 43296
rect 42668 43256 42674 43268
rect 27433 43231 27491 43237
rect 27433 43197 27445 43231
rect 27479 43228 27491 43231
rect 27479 43200 28396 43228
rect 27479 43197 27491 43200
rect 27433 43191 27491 43197
rect 25792 43132 26740 43160
rect 25130 43092 25136 43104
rect 23584 43064 25136 43092
rect 25130 43052 25136 43064
rect 25188 43052 25194 43104
rect 25314 43052 25320 43104
rect 25372 43092 25378 43104
rect 25792 43092 25820 43132
rect 27246 43120 27252 43172
rect 27304 43160 27310 43172
rect 27893 43163 27951 43169
rect 27893 43160 27905 43163
rect 27304 43132 27905 43160
rect 27304 43120 27310 43132
rect 27893 43129 27905 43132
rect 27939 43129 27951 43163
rect 28368 43160 28396 43200
rect 28442 43188 28448 43240
rect 28500 43188 28506 43240
rect 28718 43188 28724 43240
rect 28776 43228 28782 43240
rect 28813 43231 28871 43237
rect 28813 43228 28825 43231
rect 28776 43200 28825 43228
rect 28776 43188 28782 43200
rect 28813 43197 28825 43200
rect 28859 43197 28871 43231
rect 28813 43191 28871 43197
rect 29362 43188 29368 43240
rect 29420 43188 29426 43240
rect 30558 43188 30564 43240
rect 30616 43228 30622 43240
rect 30727 43231 30785 43237
rect 30727 43228 30739 43231
rect 30616 43200 30739 43228
rect 30616 43188 30622 43200
rect 30727 43197 30739 43200
rect 30773 43197 30785 43231
rect 30727 43191 30785 43197
rect 31202 43188 31208 43240
rect 31260 43188 31266 43240
rect 31570 43188 31576 43240
rect 31628 43188 31634 43240
rect 34606 43188 34612 43240
rect 34664 43228 34670 43240
rect 34701 43231 34759 43237
rect 34701 43228 34713 43231
rect 34664 43200 34713 43228
rect 34664 43188 34670 43200
rect 34701 43197 34713 43200
rect 34747 43197 34759 43231
rect 38948 43228 38976 43256
rect 39758 43228 39764 43240
rect 38948 43200 39764 43228
rect 34701 43191 34759 43197
rect 39758 43188 39764 43200
rect 39816 43228 39822 43240
rect 39853 43231 39911 43237
rect 39853 43228 39865 43231
rect 39816 43200 39865 43228
rect 39816 43188 39822 43200
rect 39853 43197 39865 43200
rect 39899 43197 39911 43231
rect 39853 43191 39911 43197
rect 40862 43188 40868 43240
rect 40920 43188 40926 43240
rect 42886 43228 42892 43240
rect 42366 43200 42892 43228
rect 42886 43188 42892 43200
rect 42944 43188 42950 43240
rect 43180 43228 43208 43268
rect 43257 43265 43269 43299
rect 43303 43265 43315 43299
rect 43257 43259 43315 43265
rect 43349 43299 43407 43305
rect 43349 43265 43361 43299
rect 43395 43265 43407 43299
rect 43349 43259 43407 43265
rect 45005 43299 45063 43305
rect 45005 43265 45017 43299
rect 45051 43265 45063 43299
rect 45005 43259 45063 43265
rect 45833 43299 45891 43305
rect 45833 43265 45845 43299
rect 45879 43296 45891 43299
rect 47210 43296 47216 43308
rect 45879 43268 47216 43296
rect 45879 43265 45891 43268
rect 45833 43259 45891 43265
rect 43364 43228 43392 43259
rect 43180 43200 43392 43228
rect 43717 43231 43775 43237
rect 43717 43197 43729 43231
rect 43763 43228 43775 43231
rect 43898 43228 43904 43240
rect 43763 43200 43904 43228
rect 43763 43197 43775 43200
rect 43717 43191 43775 43197
rect 43898 43188 43904 43200
rect 43956 43188 43962 43240
rect 45848 43228 45876 43259
rect 47210 43256 47216 43268
rect 47268 43256 47274 43308
rect 47302 43256 47308 43308
rect 47360 43256 47366 43308
rect 47673 43299 47731 43305
rect 47673 43265 47685 43299
rect 47719 43296 47731 43299
rect 48682 43296 48688 43308
rect 47719 43268 48688 43296
rect 47719 43265 47731 43268
rect 47673 43259 47731 43265
rect 48682 43256 48688 43268
rect 48740 43256 48746 43308
rect 44192 43200 45876 43228
rect 47581 43231 47639 43237
rect 28626 43160 28632 43172
rect 28368 43132 28632 43160
rect 27893 43123 27951 43129
rect 28626 43120 28632 43132
rect 28684 43120 28690 43172
rect 30190 43120 30196 43172
rect 30248 43160 30254 43172
rect 31386 43160 31392 43172
rect 30248 43132 31392 43160
rect 30248 43120 30254 43132
rect 31386 43120 31392 43132
rect 31444 43120 31450 43172
rect 33226 43120 33232 43172
rect 33284 43160 33290 43172
rect 33686 43160 33692 43172
rect 33284 43132 33692 43160
rect 33284 43120 33290 43132
rect 33686 43120 33692 43132
rect 33744 43120 33750 43172
rect 34054 43120 34060 43172
rect 34112 43160 34118 43172
rect 34112 43132 35112 43160
rect 34112 43120 34118 43132
rect 25372 43064 25820 43092
rect 25961 43095 26019 43101
rect 25372 43052 25378 43064
rect 25961 43061 25973 43095
rect 26007 43092 26019 43095
rect 26142 43092 26148 43104
rect 26007 43064 26148 43092
rect 26007 43061 26019 43064
rect 25961 43055 26019 43061
rect 26142 43052 26148 43064
rect 26200 43052 26206 43104
rect 26510 43052 26516 43104
rect 26568 43052 26574 43104
rect 27065 43095 27123 43101
rect 27065 43061 27077 43095
rect 27111 43092 27123 43095
rect 27338 43092 27344 43104
rect 27111 43064 27344 43092
rect 27111 43061 27123 43064
rect 27065 43055 27123 43061
rect 27338 43052 27344 43064
rect 27396 43052 27402 43104
rect 27430 43052 27436 43104
rect 27488 43092 27494 43104
rect 29086 43092 29092 43104
rect 27488 43064 29092 43092
rect 27488 43052 27494 43064
rect 29086 43052 29092 43064
rect 29144 43052 29150 43104
rect 29457 43095 29515 43101
rect 29457 43061 29469 43095
rect 29503 43092 29515 43095
rect 29730 43092 29736 43104
rect 29503 43064 29736 43092
rect 29503 43061 29515 43064
rect 29457 43055 29515 43061
rect 29730 43052 29736 43064
rect 29788 43052 29794 43104
rect 30282 43052 30288 43104
rect 30340 43052 30346 43104
rect 30558 43052 30564 43104
rect 30616 43092 30622 43104
rect 30837 43095 30895 43101
rect 30837 43092 30849 43095
rect 30616 43064 30849 43092
rect 30616 43052 30622 43064
rect 30837 43061 30849 43064
rect 30883 43061 30895 43095
rect 30837 43055 30895 43061
rect 32214 43052 32220 43104
rect 32272 43092 32278 43104
rect 34330 43092 34336 43104
rect 32272 43064 34336 43092
rect 32272 43052 32278 43064
rect 34330 43052 34336 43064
rect 34388 43052 34394 43104
rect 35084 43092 35112 43132
rect 35158 43120 35164 43172
rect 35216 43120 35222 43172
rect 38746 43160 38752 43172
rect 35268 43132 35650 43160
rect 38686 43132 38752 43160
rect 35268 43092 35296 43132
rect 38746 43120 38752 43132
rect 38804 43120 38810 43172
rect 40402 43120 40408 43172
rect 40460 43120 40466 43172
rect 41233 43163 41291 43169
rect 41233 43129 41245 43163
rect 41279 43160 41291 43163
rect 41506 43160 41512 43172
rect 41279 43132 41512 43160
rect 41279 43129 41291 43132
rect 41233 43123 41291 43129
rect 41506 43120 41512 43132
rect 41564 43120 41570 43172
rect 43165 43163 43223 43169
rect 43165 43160 43177 43163
rect 42536 43132 43177 43160
rect 35084 43064 35296 43092
rect 39942 43052 39948 43104
rect 40000 43092 40006 43104
rect 40681 43095 40739 43101
rect 40681 43092 40693 43095
rect 40000 43064 40693 43092
rect 40000 43052 40006 43064
rect 40681 43061 40693 43064
rect 40727 43061 40739 43095
rect 40681 43055 40739 43061
rect 41046 43052 41052 43104
rect 41104 43092 41110 43104
rect 42536 43092 42564 43132
rect 43165 43129 43177 43132
rect 43211 43129 43223 43163
rect 44192 43160 44220 43200
rect 47581 43197 47593 43231
rect 47627 43197 47639 43231
rect 47581 43191 47639 43197
rect 49421 43231 49479 43237
rect 49421 43197 49433 43231
rect 49467 43228 49479 43231
rect 49970 43228 49976 43240
rect 49467 43200 49976 43228
rect 49467 43197 49479 43200
rect 49421 43191 49479 43197
rect 43165 43123 43223 43129
rect 43364 43132 44220 43160
rect 44269 43163 44327 43169
rect 41104 43064 42564 43092
rect 41104 43052 41110 43064
rect 43070 43052 43076 43104
rect 43128 43092 43134 43104
rect 43364 43092 43392 43132
rect 44269 43129 44281 43163
rect 44315 43160 44327 43163
rect 44821 43163 44879 43169
rect 44821 43160 44833 43163
rect 44315 43132 44833 43160
rect 44315 43129 44327 43132
rect 44269 43123 44327 43129
rect 44821 43129 44833 43132
rect 44867 43129 44879 43163
rect 44821 43123 44879 43129
rect 46014 43120 46020 43172
rect 46072 43160 46078 43172
rect 46072 43132 46138 43160
rect 46072 43120 46078 43132
rect 47394 43120 47400 43172
rect 47452 43160 47458 43172
rect 47596 43160 47624 43191
rect 49970 43188 49976 43200
rect 50028 43188 50034 43240
rect 51718 43188 51724 43240
rect 51776 43228 51782 43240
rect 51813 43231 51871 43237
rect 51813 43228 51825 43231
rect 51776 43200 51825 43228
rect 51776 43188 51782 43200
rect 51813 43197 51825 43200
rect 51859 43197 51871 43231
rect 51813 43191 51871 43197
rect 47452 43132 47624 43160
rect 47452 43120 47458 43132
rect 48130 43120 48136 43172
rect 48188 43120 48194 43172
rect 49142 43120 49148 43172
rect 49200 43120 49206 43172
rect 52362 43120 52368 43172
rect 52420 43120 52426 43172
rect 43128 43064 43392 43092
rect 43128 43052 43134 43064
rect 43438 43052 43444 43104
rect 43496 43092 43502 43104
rect 44453 43095 44511 43101
rect 44453 43092 44465 43095
rect 43496 43064 44465 43092
rect 43496 43052 43502 43064
rect 44453 43061 44465 43064
rect 44499 43061 44511 43095
rect 44453 43055 44511 43061
rect 44910 43052 44916 43104
rect 44968 43052 44974 43104
rect 51261 43095 51319 43101
rect 51261 43061 51273 43095
rect 51307 43092 51319 43095
rect 51534 43092 51540 43104
rect 51307 43064 51540 43092
rect 51307 43061 51319 43064
rect 51261 43055 51319 43061
rect 51534 43052 51540 43064
rect 51592 43052 51598 43104
rect 51810 43052 51816 43104
rect 51868 43092 51874 43104
rect 52089 43095 52147 43101
rect 52089 43092 52101 43095
rect 51868 43064 52101 43092
rect 51868 43052 51874 43064
rect 52089 43061 52101 43064
rect 52135 43061 52147 43095
rect 52089 43055 52147 43061
rect 552 43002 66424 43024
rect 552 42950 2918 43002
rect 2970 42950 2982 43002
rect 3034 42950 3046 43002
rect 3098 42950 3110 43002
rect 3162 42950 3174 43002
rect 3226 42950 51918 43002
rect 51970 42950 51982 43002
rect 52034 42950 52046 43002
rect 52098 42950 52110 43002
rect 52162 42950 52174 43002
rect 52226 42950 66424 43002
rect 552 42928 66424 42950
rect 11698 42848 11704 42900
rect 11756 42888 11762 42900
rect 12069 42891 12127 42897
rect 12069 42888 12081 42891
rect 11756 42860 12081 42888
rect 11756 42848 11762 42860
rect 12069 42857 12081 42860
rect 12115 42857 12127 42891
rect 12069 42851 12127 42857
rect 12250 42848 12256 42900
rect 12308 42888 12314 42900
rect 12437 42891 12495 42897
rect 12437 42888 12449 42891
rect 12308 42860 12449 42888
rect 12308 42848 12314 42860
rect 12437 42857 12449 42860
rect 12483 42857 12495 42891
rect 12437 42851 12495 42857
rect 12526 42848 12532 42900
rect 12584 42888 12590 42900
rect 12897 42891 12955 42897
rect 12897 42888 12909 42891
rect 12584 42860 12909 42888
rect 12584 42848 12590 42860
rect 12897 42857 12909 42860
rect 12943 42857 12955 42891
rect 12897 42851 12955 42857
rect 13357 42891 13415 42897
rect 13357 42857 13369 42891
rect 13403 42888 13415 42891
rect 13998 42888 14004 42900
rect 13403 42860 14004 42888
rect 13403 42857 13415 42860
rect 13357 42851 13415 42857
rect 13998 42848 14004 42860
rect 14056 42848 14062 42900
rect 14093 42891 14151 42897
rect 14093 42857 14105 42891
rect 14139 42888 14151 42891
rect 14366 42888 14372 42900
rect 14139 42860 14372 42888
rect 14139 42857 14151 42860
rect 14093 42851 14151 42857
rect 14366 42848 14372 42860
rect 14424 42848 14430 42900
rect 14734 42848 14740 42900
rect 14792 42888 14798 42900
rect 16206 42888 16212 42900
rect 14792 42860 16212 42888
rect 14792 42848 14798 42860
rect 16206 42848 16212 42860
rect 16264 42888 16270 42900
rect 19518 42888 19524 42900
rect 16264 42860 19524 42888
rect 16264 42848 16270 42860
rect 14182 42780 14188 42832
rect 14240 42820 14246 42832
rect 16666 42820 16672 42832
rect 14240 42792 14780 42820
rect 14240 42780 14246 42792
rect 12529 42755 12587 42761
rect 12529 42721 12541 42755
rect 12575 42752 12587 42755
rect 13170 42752 13176 42764
rect 12575 42724 13176 42752
rect 12575 42721 12587 42724
rect 12529 42715 12587 42721
rect 13170 42712 13176 42724
rect 13228 42752 13234 42764
rect 13265 42755 13323 42761
rect 13265 42752 13277 42755
rect 13228 42724 13277 42752
rect 13228 42712 13234 42724
rect 13265 42721 13277 42724
rect 13311 42752 13323 42755
rect 14550 42752 14556 42764
rect 13311 42724 14556 42752
rect 13311 42721 13323 42724
rect 13265 42715 13323 42721
rect 14550 42712 14556 42724
rect 14608 42712 14614 42764
rect 14752 42761 14780 42792
rect 16040 42792 16672 42820
rect 14737 42755 14795 42761
rect 14737 42721 14749 42755
rect 14783 42752 14795 42755
rect 15010 42752 15016 42764
rect 14783 42724 15016 42752
rect 14783 42721 14795 42724
rect 14737 42715 14795 42721
rect 15010 42712 15016 42724
rect 15068 42712 15074 42764
rect 15197 42755 15255 42761
rect 15197 42721 15209 42755
rect 15243 42752 15255 42755
rect 16040 42752 16068 42792
rect 16666 42780 16672 42792
rect 16724 42780 16730 42832
rect 16942 42780 16948 42832
rect 17000 42780 17006 42832
rect 15243 42724 16068 42752
rect 15243 42721 15255 42724
rect 15197 42715 15255 42721
rect 16114 42712 16120 42764
rect 16172 42712 16178 42764
rect 18432 42761 18460 42860
rect 19518 42848 19524 42860
rect 19576 42888 19582 42900
rect 19978 42888 19984 42900
rect 19576 42860 19984 42888
rect 19576 42848 19582 42860
rect 19978 42848 19984 42860
rect 20036 42848 20042 42900
rect 20254 42848 20260 42900
rect 20312 42848 20318 42900
rect 20717 42891 20775 42897
rect 20717 42857 20729 42891
rect 20763 42888 20775 42891
rect 20806 42888 20812 42900
rect 20763 42860 20812 42888
rect 20763 42857 20775 42860
rect 20717 42851 20775 42857
rect 20162 42820 20168 42832
rect 19918 42792 20168 42820
rect 20162 42780 20168 42792
rect 20220 42780 20226 42832
rect 20732 42820 20760 42851
rect 20806 42848 20812 42860
rect 20864 42848 20870 42900
rect 22005 42891 22063 42897
rect 22005 42857 22017 42891
rect 22051 42888 22063 42891
rect 22554 42888 22560 42900
rect 22051 42860 22560 42888
rect 22051 42857 22063 42860
rect 22005 42851 22063 42857
rect 22554 42848 22560 42860
rect 22612 42848 22618 42900
rect 22738 42848 22744 42900
rect 22796 42848 22802 42900
rect 24210 42848 24216 42900
rect 24268 42888 24274 42900
rect 24857 42891 24915 42897
rect 24857 42888 24869 42891
rect 24268 42860 24869 42888
rect 24268 42848 24274 42860
rect 24857 42857 24869 42860
rect 24903 42888 24915 42891
rect 25406 42888 25412 42900
rect 24903 42860 25412 42888
rect 24903 42857 24915 42860
rect 24857 42851 24915 42857
rect 25406 42848 25412 42860
rect 25464 42848 25470 42900
rect 25777 42891 25835 42897
rect 25777 42857 25789 42891
rect 25823 42888 25835 42891
rect 26142 42888 26148 42900
rect 25823 42860 26148 42888
rect 25823 42857 25835 42860
rect 25777 42851 25835 42857
rect 26142 42848 26148 42860
rect 26200 42848 26206 42900
rect 26237 42891 26295 42897
rect 26237 42857 26249 42891
rect 26283 42888 26295 42891
rect 26510 42888 26516 42900
rect 26283 42860 26516 42888
rect 26283 42857 26295 42860
rect 26237 42851 26295 42857
rect 26510 42848 26516 42860
rect 26568 42848 26574 42900
rect 27706 42848 27712 42900
rect 27764 42888 27770 42900
rect 38562 42888 38568 42900
rect 27764 42860 38568 42888
rect 27764 42848 27770 42860
rect 38562 42848 38568 42860
rect 38620 42848 38626 42900
rect 38654 42848 38660 42900
rect 38712 42848 38718 42900
rect 39022 42848 39028 42900
rect 39080 42848 39086 42900
rect 39117 42891 39175 42897
rect 39117 42857 39129 42891
rect 39163 42888 39175 42891
rect 39298 42888 39304 42900
rect 39163 42860 39304 42888
rect 39163 42857 39175 42860
rect 39117 42851 39175 42857
rect 39298 42848 39304 42860
rect 39356 42848 39362 42900
rect 40313 42891 40371 42897
rect 40313 42857 40325 42891
rect 40359 42888 40371 42891
rect 40402 42888 40408 42900
rect 40359 42860 40408 42888
rect 40359 42857 40371 42860
rect 40313 42851 40371 42857
rect 40402 42848 40408 42860
rect 40460 42888 40466 42900
rect 40770 42888 40776 42900
rect 40460 42860 40776 42888
rect 40460 42848 40466 42860
rect 40770 42848 40776 42860
rect 40828 42848 40834 42900
rect 41046 42848 41052 42900
rect 41104 42848 41110 42900
rect 41414 42848 41420 42900
rect 41472 42848 41478 42900
rect 43806 42848 43812 42900
rect 43864 42888 43870 42900
rect 44361 42891 44419 42897
rect 44361 42888 44373 42891
rect 43864 42860 44373 42888
rect 43864 42848 43870 42860
rect 44361 42857 44373 42860
rect 44407 42857 44419 42891
rect 44361 42851 44419 42857
rect 44729 42891 44787 42897
rect 44729 42857 44741 42891
rect 44775 42888 44787 42891
rect 44910 42888 44916 42900
rect 44775 42860 44916 42888
rect 44775 42857 44787 42860
rect 44729 42851 44787 42857
rect 44910 42848 44916 42860
rect 44968 42848 44974 42900
rect 46014 42848 46020 42900
rect 46072 42888 46078 42900
rect 46569 42891 46627 42897
rect 46569 42888 46581 42891
rect 46072 42860 46581 42888
rect 46072 42848 46078 42860
rect 46569 42857 46581 42860
rect 46615 42857 46627 42891
rect 46569 42851 46627 42857
rect 46934 42848 46940 42900
rect 46992 42888 46998 42900
rect 47029 42891 47087 42897
rect 47029 42888 47041 42891
rect 46992 42860 47041 42888
rect 46992 42848 46998 42860
rect 47029 42857 47041 42860
rect 47075 42857 47087 42891
rect 47029 42851 47087 42857
rect 47210 42848 47216 42900
rect 47268 42888 47274 42900
rect 47397 42891 47455 42897
rect 47397 42888 47409 42891
rect 47268 42860 47409 42888
rect 47268 42848 47274 42860
rect 47397 42857 47409 42860
rect 47443 42857 47455 42891
rect 47397 42851 47455 42857
rect 48593 42891 48651 42897
rect 48593 42857 48605 42891
rect 48639 42888 48651 42891
rect 48682 42888 48688 42900
rect 48639 42860 48688 42888
rect 48639 42857 48651 42860
rect 48593 42851 48651 42857
rect 48682 42848 48688 42860
rect 48740 42848 48746 42900
rect 49053 42891 49111 42897
rect 49053 42857 49065 42891
rect 49099 42888 49111 42891
rect 49142 42888 49148 42900
rect 49099 42860 49148 42888
rect 49099 42857 49111 42860
rect 49053 42851 49111 42857
rect 49142 42848 49148 42860
rect 49200 42848 49206 42900
rect 49418 42848 49424 42900
rect 49476 42848 49482 42900
rect 20548 42792 20760 42820
rect 21637 42823 21695 42829
rect 18417 42755 18475 42761
rect 18417 42721 18429 42755
rect 18463 42721 18475 42755
rect 18417 42715 18475 42721
rect 12713 42687 12771 42693
rect 12713 42653 12725 42687
rect 12759 42684 12771 42687
rect 13078 42684 13084 42696
rect 12759 42656 13084 42684
rect 12759 42653 12771 42656
rect 12713 42647 12771 42653
rect 13078 42644 13084 42656
rect 13136 42644 13142 42696
rect 13538 42644 13544 42696
rect 13596 42644 13602 42696
rect 13998 42644 14004 42696
rect 14056 42684 14062 42696
rect 14185 42687 14243 42693
rect 14185 42684 14197 42687
rect 14056 42656 14197 42684
rect 14056 42644 14062 42656
rect 14185 42653 14197 42656
rect 14231 42653 14243 42687
rect 14185 42647 14243 42653
rect 14369 42687 14427 42693
rect 14369 42653 14381 42687
rect 14415 42684 14427 42687
rect 14642 42684 14648 42696
rect 14415 42656 14648 42684
rect 14415 42653 14427 42656
rect 14369 42647 14427 42653
rect 14642 42644 14648 42656
rect 14700 42644 14706 42696
rect 15378 42644 15384 42696
rect 15436 42644 15442 42696
rect 16393 42687 16451 42693
rect 16393 42653 16405 42687
rect 16439 42684 16451 42687
rect 16758 42684 16764 42696
rect 16439 42656 16764 42684
rect 16439 42653 16451 42656
rect 16393 42647 16451 42653
rect 16758 42644 16764 42656
rect 16816 42644 16822 42696
rect 18693 42687 18751 42693
rect 18693 42653 18705 42687
rect 18739 42684 18751 42687
rect 19426 42684 19432 42696
rect 18739 42656 19432 42684
rect 18739 42653 18751 42656
rect 18693 42647 18751 42653
rect 19426 42644 19432 42656
rect 19484 42644 19490 42696
rect 20165 42687 20223 42693
rect 20165 42653 20177 42687
rect 20211 42684 20223 42687
rect 20548 42684 20576 42792
rect 21637 42789 21649 42823
rect 21683 42820 21695 42823
rect 22094 42820 22100 42832
rect 21683 42792 22100 42820
rect 21683 42789 21695 42792
rect 21637 42783 21695 42789
rect 22094 42780 22100 42792
rect 22152 42780 22158 42832
rect 24946 42820 24952 42832
rect 24610 42792 24952 42820
rect 24946 42780 24952 42792
rect 25004 42780 25010 42832
rect 27246 42780 27252 42832
rect 27304 42780 27310 42832
rect 27338 42780 27344 42832
rect 27396 42780 27402 42832
rect 28077 42823 28135 42829
rect 28077 42789 28089 42823
rect 28123 42820 28135 42823
rect 28994 42820 29000 42832
rect 28123 42792 29000 42820
rect 28123 42789 28135 42792
rect 28077 42783 28135 42789
rect 28994 42780 29000 42792
rect 29052 42780 29058 42832
rect 29365 42823 29423 42829
rect 29365 42789 29377 42823
rect 29411 42820 29423 42823
rect 30190 42820 30196 42832
rect 29411 42792 30196 42820
rect 29411 42789 29423 42792
rect 29365 42783 29423 42789
rect 30190 42780 30196 42792
rect 30248 42780 30254 42832
rect 30374 42780 30380 42832
rect 30432 42820 30438 42832
rect 30561 42823 30619 42829
rect 30561 42820 30573 42823
rect 30432 42792 30573 42820
rect 30432 42780 30438 42792
rect 30561 42789 30573 42792
rect 30607 42789 30619 42823
rect 30561 42783 30619 42789
rect 32398 42780 32404 42832
rect 32456 42780 32462 42832
rect 33686 42820 33692 42832
rect 33626 42792 33692 42820
rect 33686 42780 33692 42792
rect 33744 42820 33750 42832
rect 34146 42820 34152 42832
rect 33744 42792 34152 42820
rect 33744 42780 33750 42792
rect 34146 42780 34152 42792
rect 34204 42780 34210 42832
rect 34330 42780 34336 42832
rect 34388 42780 34394 42832
rect 35345 42823 35403 42829
rect 35345 42789 35357 42823
rect 35391 42820 35403 42823
rect 35526 42820 35532 42832
rect 35391 42792 35532 42820
rect 35391 42789 35403 42792
rect 35345 42783 35403 42789
rect 35526 42780 35532 42792
rect 35584 42780 35590 42832
rect 37369 42823 37427 42829
rect 37369 42820 37381 42823
rect 36832 42792 37381 42820
rect 36832 42764 36860 42792
rect 37369 42789 37381 42792
rect 37415 42789 37427 42823
rect 37369 42783 37427 42789
rect 38197 42823 38255 42829
rect 38197 42789 38209 42823
rect 38243 42820 38255 42823
rect 39485 42823 39543 42829
rect 39485 42820 39497 42823
rect 38243 42792 39497 42820
rect 38243 42789 38255 42792
rect 38197 42783 38255 42789
rect 39485 42789 39497 42792
rect 39531 42789 39543 42823
rect 39485 42783 39543 42789
rect 39942 42780 39948 42832
rect 40000 42820 40006 42832
rect 42886 42820 42892 42832
rect 40000 42792 42892 42820
rect 40000 42780 40006 42792
rect 42886 42780 42892 42792
rect 42944 42780 42950 42832
rect 51810 42820 51816 42832
rect 51474 42792 51816 42820
rect 51810 42780 51816 42792
rect 51868 42780 51874 42832
rect 20625 42755 20683 42761
rect 20625 42721 20637 42755
rect 20671 42752 20683 42755
rect 20898 42752 20904 42764
rect 20671 42724 20904 42752
rect 20671 42721 20683 42724
rect 20625 42715 20683 42721
rect 20898 42712 20904 42724
rect 20956 42712 20962 42764
rect 22370 42712 22376 42764
rect 22428 42752 22434 42764
rect 22649 42755 22707 42761
rect 22649 42752 22661 42755
rect 22428 42724 22661 42752
rect 22428 42712 22434 42724
rect 22649 42721 22661 42724
rect 22695 42721 22707 42755
rect 22649 42715 22707 42721
rect 25866 42712 25872 42764
rect 25924 42712 25930 42764
rect 26418 42712 26424 42764
rect 26476 42712 26482 42764
rect 27540 42724 28396 42752
rect 20211 42656 20576 42684
rect 20809 42687 20867 42693
rect 20211 42653 20223 42656
rect 20165 42647 20223 42653
rect 20809 42653 20821 42687
rect 20855 42653 20867 42687
rect 20809 42647 20867 42653
rect 13725 42619 13783 42625
rect 13725 42585 13737 42619
rect 13771 42616 13783 42619
rect 13814 42616 13820 42628
rect 13771 42588 13820 42616
rect 13771 42585 13783 42588
rect 13725 42579 13783 42585
rect 13814 42576 13820 42588
rect 13872 42576 13878 42628
rect 15010 42576 15016 42628
rect 15068 42576 15074 42628
rect 20824 42616 20852 42647
rect 21450 42644 21456 42696
rect 21508 42644 21514 42696
rect 21545 42687 21603 42693
rect 21545 42653 21557 42687
rect 21591 42684 21603 42687
rect 21591 42656 22094 42684
rect 21591 42653 21603 42656
rect 21545 42647 21603 42653
rect 20732 42588 20852 42616
rect 22066 42616 22094 42656
rect 22554 42644 22560 42696
rect 22612 42684 22618 42696
rect 22830 42684 22836 42696
rect 22612 42656 22836 42684
rect 22612 42644 22618 42656
rect 22830 42644 22836 42656
rect 22888 42644 22894 42696
rect 23109 42687 23167 42693
rect 23109 42653 23121 42687
rect 23155 42653 23167 42687
rect 23109 42647 23167 42653
rect 22281 42619 22339 42625
rect 22281 42616 22293 42619
rect 22066 42588 22293 42616
rect 14274 42508 14280 42560
rect 14332 42548 14338 42560
rect 14645 42551 14703 42557
rect 14645 42548 14657 42551
rect 14332 42520 14657 42548
rect 14332 42508 14338 42520
rect 14645 42517 14657 42520
rect 14691 42517 14703 42551
rect 14645 42511 14703 42517
rect 15933 42551 15991 42557
rect 15933 42517 15945 42551
rect 15979 42548 15991 42551
rect 17126 42548 17132 42560
rect 15979 42520 17132 42548
rect 15979 42517 15991 42520
rect 15933 42511 15991 42517
rect 17126 42508 17132 42520
rect 17184 42508 17190 42560
rect 17865 42551 17923 42557
rect 17865 42517 17877 42551
rect 17911 42548 17923 42551
rect 17954 42548 17960 42560
rect 17911 42520 17960 42548
rect 17911 42517 17923 42520
rect 17865 42511 17923 42517
rect 17954 42508 17960 42520
rect 18012 42508 18018 42560
rect 19242 42508 19248 42560
rect 19300 42548 19306 42560
rect 20732 42548 20760 42588
rect 22281 42585 22293 42588
rect 22327 42585 22339 42619
rect 22281 42579 22339 42585
rect 20806 42548 20812 42560
rect 19300 42520 20812 42548
rect 19300 42508 19306 42520
rect 20806 42508 20812 42520
rect 20864 42508 20870 42560
rect 22189 42551 22247 42557
rect 22189 42517 22201 42551
rect 22235 42548 22247 42551
rect 22370 42548 22376 42560
rect 22235 42520 22376 42548
rect 22235 42517 22247 42520
rect 22189 42511 22247 42517
rect 22370 42508 22376 42520
rect 22428 42508 22434 42560
rect 23124 42548 23152 42647
rect 23382 42644 23388 42696
rect 23440 42644 23446 42696
rect 25685 42687 25743 42693
rect 25685 42653 25697 42687
rect 25731 42684 25743 42687
rect 26050 42684 26056 42696
rect 25731 42656 26056 42684
rect 25731 42653 25743 42656
rect 25685 42647 25743 42653
rect 26050 42644 26056 42656
rect 26108 42644 26114 42696
rect 27540 42693 27568 42724
rect 28368 42696 28396 42724
rect 28810 42712 28816 42764
rect 28868 42712 28874 42764
rect 29273 42755 29331 42761
rect 29273 42752 29285 42755
rect 28920 42724 29285 42752
rect 27525 42687 27583 42693
rect 26344 42656 27384 42684
rect 24670 42576 24676 42628
rect 24728 42616 24734 42628
rect 26344 42616 26372 42656
rect 24728 42588 26372 42616
rect 24728 42576 24734 42588
rect 26602 42576 26608 42628
rect 26660 42576 26666 42628
rect 23474 42548 23480 42560
rect 23124 42520 23480 42548
rect 23474 42508 23480 42520
rect 23532 42508 23538 42560
rect 26694 42508 26700 42560
rect 26752 42548 26758 42560
rect 26881 42551 26939 42557
rect 26881 42548 26893 42551
rect 26752 42520 26893 42548
rect 26752 42508 26758 42520
rect 26881 42517 26893 42520
rect 26927 42517 26939 42551
rect 27356 42548 27384 42656
rect 27525 42653 27537 42687
rect 27571 42653 27583 42687
rect 27525 42647 27583 42653
rect 27614 42644 27620 42696
rect 27672 42684 27678 42696
rect 27672 42656 27752 42684
rect 27672 42644 27678 42656
rect 27724 42625 27752 42656
rect 28166 42644 28172 42696
rect 28224 42644 28230 42696
rect 28350 42644 28356 42696
rect 28408 42644 28414 42696
rect 28626 42644 28632 42696
rect 28684 42684 28690 42696
rect 28920 42684 28948 42724
rect 29273 42721 29285 42724
rect 29319 42721 29331 42755
rect 29273 42715 29331 42721
rect 30466 42712 30472 42764
rect 30524 42752 30530 42764
rect 30653 42755 30711 42761
rect 30653 42752 30665 42755
rect 30524 42724 30665 42752
rect 30524 42712 30530 42724
rect 30653 42721 30665 42724
rect 30699 42721 30711 42755
rect 30653 42715 30711 42721
rect 35066 42712 35072 42764
rect 35124 42752 35130 42764
rect 35437 42755 35495 42761
rect 35437 42752 35449 42755
rect 35124 42724 35449 42752
rect 35124 42712 35130 42724
rect 35437 42721 35449 42724
rect 35483 42721 35495 42755
rect 35437 42715 35495 42721
rect 36541 42755 36599 42761
rect 36541 42721 36553 42755
rect 36587 42752 36599 42755
rect 36630 42752 36636 42764
rect 36587 42724 36636 42752
rect 36587 42721 36599 42724
rect 36541 42715 36599 42721
rect 36630 42712 36636 42724
rect 36688 42712 36694 42764
rect 36814 42712 36820 42764
rect 36872 42712 36878 42764
rect 37274 42712 37280 42764
rect 37332 42712 37338 42764
rect 38289 42755 38347 42761
rect 38289 42721 38301 42755
rect 38335 42752 38347 42755
rect 39114 42752 39120 42764
rect 38335 42724 39120 42752
rect 38335 42721 38347 42724
rect 38289 42715 38347 42721
rect 39114 42712 39120 42724
rect 39172 42712 39178 42764
rect 40494 42712 40500 42764
rect 40552 42712 40558 42764
rect 41322 42712 41328 42764
rect 41380 42752 41386 42764
rect 42153 42755 42211 42761
rect 42153 42752 42165 42755
rect 41380 42724 42165 42752
rect 41380 42712 41386 42724
rect 42153 42721 42165 42724
rect 42199 42721 42211 42755
rect 42153 42715 42211 42721
rect 43714 42712 43720 42764
rect 43772 42752 43778 42764
rect 44913 42755 44971 42761
rect 44913 42752 44925 42755
rect 43772 42724 44925 42752
rect 43772 42712 43778 42724
rect 44913 42721 44925 42724
rect 44959 42721 44971 42755
rect 44913 42715 44971 42721
rect 46477 42755 46535 42761
rect 46477 42721 46489 42755
rect 46523 42752 46535 42755
rect 46566 42752 46572 42764
rect 46523 42724 46572 42752
rect 46523 42721 46535 42724
rect 46477 42715 46535 42721
rect 46566 42712 46572 42724
rect 46624 42752 46630 42764
rect 48130 42752 48136 42764
rect 46624 42724 48136 42752
rect 46624 42712 46630 42724
rect 48130 42712 48136 42724
rect 48188 42712 48194 42764
rect 48222 42712 48228 42764
rect 48280 42752 48286 42764
rect 48280 42724 49648 42752
rect 48280 42712 48286 42724
rect 28684 42656 28948 42684
rect 28684 42644 28690 42656
rect 29086 42644 29092 42696
rect 29144 42684 29150 42696
rect 30745 42687 30803 42693
rect 30745 42684 30757 42687
rect 29144 42656 30757 42684
rect 29144 42644 29150 42656
rect 30745 42653 30757 42656
rect 30791 42653 30803 42687
rect 30745 42647 30803 42653
rect 32122 42644 32128 42696
rect 32180 42644 32186 42696
rect 33686 42644 33692 42696
rect 33744 42684 33750 42696
rect 34425 42687 34483 42693
rect 34425 42684 34437 42687
rect 33744 42656 34437 42684
rect 33744 42644 33750 42656
rect 34425 42653 34437 42656
rect 34471 42653 34483 42687
rect 34425 42647 34483 42653
rect 34514 42644 34520 42696
rect 34572 42644 34578 42696
rect 34974 42644 34980 42696
rect 35032 42684 35038 42696
rect 35161 42687 35219 42693
rect 35161 42684 35173 42687
rect 35032 42656 35173 42684
rect 35032 42644 35038 42656
rect 35161 42653 35173 42656
rect 35207 42653 35219 42687
rect 37185 42687 37243 42693
rect 37185 42684 37197 42687
rect 35161 42647 35219 42653
rect 35866 42656 37197 42684
rect 27709 42619 27767 42625
rect 27709 42585 27721 42619
rect 27755 42585 27767 42619
rect 27709 42579 27767 42585
rect 27798 42576 27804 42628
rect 27856 42616 27862 42628
rect 29178 42616 29184 42628
rect 27856 42588 29184 42616
rect 27856 42576 27862 42588
rect 29178 42576 29184 42588
rect 29236 42576 29242 42628
rect 29730 42576 29736 42628
rect 29788 42576 29794 42628
rect 30193 42619 30251 42625
rect 30193 42585 30205 42619
rect 30239 42616 30251 42619
rect 30282 42616 30288 42628
rect 30239 42588 30288 42616
rect 30239 42585 30251 42588
rect 30193 42579 30251 42585
rect 30282 42576 30288 42588
rect 30340 42576 30346 42628
rect 33410 42576 33416 42628
rect 33468 42616 33474 42628
rect 33965 42619 34023 42625
rect 33965 42616 33977 42619
rect 33468 42588 33977 42616
rect 33468 42576 33474 42588
rect 33965 42585 33977 42588
rect 34011 42585 34023 42619
rect 34532 42616 34560 42644
rect 35866 42616 35894 42656
rect 37185 42653 37197 42656
rect 37231 42684 37243 42687
rect 37550 42684 37556 42696
rect 37231 42656 37556 42684
rect 37231 42653 37243 42656
rect 37185 42647 37243 42653
rect 37550 42644 37556 42656
rect 37608 42644 37614 42696
rect 38010 42644 38016 42696
rect 38068 42684 38074 42696
rect 38378 42684 38384 42696
rect 38068 42656 38384 42684
rect 38068 42644 38074 42656
rect 38378 42644 38384 42656
rect 38436 42684 38442 42696
rect 38473 42687 38531 42693
rect 38473 42684 38485 42687
rect 38436 42656 38485 42684
rect 38436 42644 38442 42656
rect 38473 42653 38485 42656
rect 38519 42684 38531 42687
rect 39209 42687 39267 42693
rect 39209 42684 39221 42687
rect 38519 42656 39221 42684
rect 38519 42653 38531 42656
rect 38473 42647 38531 42653
rect 39209 42653 39221 42656
rect 39255 42653 39267 42687
rect 39209 42647 39267 42653
rect 34532 42588 35894 42616
rect 33965 42579 34023 42585
rect 37734 42576 37740 42628
rect 37792 42576 37798 42628
rect 39224 42616 39252 42647
rect 39298 42644 39304 42696
rect 39356 42684 39362 42696
rect 40037 42687 40095 42693
rect 40037 42684 40049 42687
rect 39356 42656 40049 42684
rect 39356 42644 39362 42656
rect 40037 42653 40049 42656
rect 40083 42653 40095 42687
rect 40037 42647 40095 42653
rect 40865 42687 40923 42693
rect 40865 42653 40877 42687
rect 40911 42653 40923 42687
rect 40865 42647 40923 42653
rect 40957 42687 41015 42693
rect 40957 42653 40969 42687
rect 41003 42684 41015 42687
rect 42058 42684 42064 42696
rect 41003 42656 42064 42684
rect 41003 42653 41015 42656
rect 40957 42647 41015 42653
rect 40880 42616 40908 42647
rect 42058 42644 42064 42656
rect 42116 42644 42122 42696
rect 42429 42687 42487 42693
rect 42429 42653 42441 42687
rect 42475 42684 42487 42687
rect 43438 42684 43444 42696
rect 42475 42656 43444 42684
rect 42475 42653 42487 42656
rect 42429 42647 42487 42653
rect 43438 42644 43444 42656
rect 43496 42644 43502 42696
rect 44174 42684 44180 42696
rect 43548 42656 44180 42684
rect 41598 42616 41604 42628
rect 39224 42588 41604 42616
rect 41598 42576 41604 42588
rect 41656 42576 41662 42628
rect 28629 42551 28687 42557
rect 28629 42548 28641 42551
rect 27356 42520 28641 42548
rect 26881 42511 26939 42517
rect 28629 42517 28641 42520
rect 28675 42548 28687 42551
rect 30098 42548 30104 42560
rect 28675 42520 30104 42548
rect 28675 42517 28687 42520
rect 28629 42511 28687 42517
rect 30098 42508 30104 42520
rect 30156 42508 30162 42560
rect 33873 42551 33931 42557
rect 33873 42517 33885 42551
rect 33919 42548 33931 42551
rect 34606 42548 34612 42560
rect 33919 42520 34612 42548
rect 33919 42517 33931 42520
rect 33873 42511 33931 42517
rect 34606 42508 34612 42520
rect 34664 42508 34670 42560
rect 34977 42551 35035 42557
rect 34977 42517 34989 42551
rect 35023 42548 35035 42551
rect 35066 42548 35072 42560
rect 35023 42520 35072 42548
rect 35023 42517 35035 42520
rect 34977 42511 35035 42517
rect 35066 42508 35072 42520
rect 35124 42508 35130 42560
rect 35710 42508 35716 42560
rect 35768 42548 35774 42560
rect 35805 42551 35863 42557
rect 35805 42548 35817 42551
rect 35768 42520 35817 42548
rect 35768 42508 35774 42520
rect 35805 42517 35817 42520
rect 35851 42517 35863 42551
rect 35805 42511 35863 42517
rect 35894 42508 35900 42560
rect 35952 42508 35958 42560
rect 37826 42508 37832 42560
rect 37884 42508 37890 42560
rect 40494 42508 40500 42560
rect 40552 42548 40558 42560
rect 42518 42548 42524 42560
rect 40552 42520 42524 42548
rect 40552 42508 40558 42520
rect 42518 42508 42524 42520
rect 42576 42508 42582 42560
rect 42610 42508 42616 42560
rect 42668 42548 42674 42560
rect 43548 42548 43576 42656
rect 44174 42644 44180 42656
rect 44232 42644 44238 42696
rect 44269 42687 44327 42693
rect 44269 42653 44281 42687
rect 44315 42653 44327 42687
rect 44269 42647 44327 42653
rect 45557 42687 45615 42693
rect 45557 42653 45569 42687
rect 45603 42684 45615 42687
rect 45646 42684 45652 42696
rect 45603 42656 45652 42684
rect 45603 42653 45615 42656
rect 45557 42647 45615 42653
rect 44284 42616 44312 42647
rect 45646 42644 45652 42656
rect 45704 42644 45710 42696
rect 46293 42687 46351 42693
rect 46293 42653 46305 42687
rect 46339 42684 46351 42687
rect 46382 42684 46388 42696
rect 46339 42656 46388 42684
rect 46339 42653 46351 42656
rect 46293 42647 46351 42653
rect 46308 42616 46336 42647
rect 46382 42644 46388 42656
rect 46440 42644 46446 42696
rect 47486 42644 47492 42696
rect 47544 42644 47550 42696
rect 47673 42687 47731 42693
rect 47673 42653 47685 42687
rect 47719 42684 47731 42687
rect 47762 42684 47768 42696
rect 47719 42656 47768 42684
rect 47719 42653 47731 42656
rect 47673 42647 47731 42653
rect 47762 42644 47768 42656
rect 47820 42644 47826 42696
rect 48682 42644 48688 42696
rect 48740 42644 48746 42696
rect 48869 42687 48927 42693
rect 48869 42653 48881 42687
rect 48915 42653 48927 42687
rect 48869 42647 48927 42653
rect 44284 42588 46336 42616
rect 47578 42576 47584 42628
rect 47636 42616 47642 42628
rect 47636 42588 48728 42616
rect 47636 42576 47642 42588
rect 42668 42520 43576 42548
rect 42668 42508 42674 42520
rect 43898 42508 43904 42560
rect 43956 42508 43962 42560
rect 44082 42508 44088 42560
rect 44140 42548 44146 42560
rect 45649 42551 45707 42557
rect 45649 42548 45661 42551
rect 44140 42520 45661 42548
rect 44140 42508 44146 42520
rect 45649 42517 45661 42520
rect 45695 42517 45707 42551
rect 45649 42511 45707 42517
rect 47670 42508 47676 42560
rect 47728 42548 47734 42560
rect 48225 42551 48283 42557
rect 48225 42548 48237 42551
rect 47728 42520 48237 42548
rect 47728 42508 47734 42520
rect 48225 42517 48237 42520
rect 48271 42517 48283 42551
rect 48700 42548 48728 42588
rect 48774 42548 48780 42560
rect 48700 42520 48780 42548
rect 48225 42511 48283 42517
rect 48774 42508 48780 42520
rect 48832 42548 48838 42560
rect 48884 42548 48912 42647
rect 49510 42644 49516 42696
rect 49568 42644 49574 42696
rect 49620 42693 49648 42724
rect 49970 42712 49976 42764
rect 50028 42712 50034 42764
rect 51626 42712 51632 42764
rect 51684 42752 51690 42764
rect 52181 42755 52239 42761
rect 52181 42752 52193 42755
rect 51684 42724 52193 42752
rect 51684 42712 51690 42724
rect 52181 42721 52193 42724
rect 52227 42752 52239 42755
rect 59998 42752 60004 42764
rect 52227 42724 60004 42752
rect 52227 42721 52239 42724
rect 52181 42715 52239 42721
rect 59998 42712 60004 42724
rect 60056 42712 60062 42764
rect 49605 42687 49663 42693
rect 49605 42653 49617 42687
rect 49651 42653 49663 42687
rect 49605 42647 49663 42653
rect 50246 42644 50252 42696
rect 50304 42644 50310 42696
rect 50338 42644 50344 42696
rect 50396 42684 50402 42696
rect 50798 42684 50804 42696
rect 50396 42656 50804 42684
rect 50396 42644 50402 42656
rect 50798 42644 50804 42656
rect 50856 42684 50862 42696
rect 54018 42684 54024 42696
rect 50856 42656 54024 42684
rect 50856 42644 50862 42656
rect 54018 42644 54024 42656
rect 54076 42644 54082 42696
rect 54110 42644 54116 42696
rect 54168 42644 54174 42696
rect 52362 42576 52368 42628
rect 52420 42616 52426 42628
rect 52420 42588 55214 42616
rect 52420 42576 52426 42588
rect 48832 42520 48912 42548
rect 48832 42508 48838 42520
rect 51718 42508 51724 42560
rect 51776 42508 51782 42560
rect 53098 42508 53104 42560
rect 53156 42548 53162 42560
rect 53561 42551 53619 42557
rect 53561 42548 53573 42551
rect 53156 42520 53573 42548
rect 53156 42508 53162 42520
rect 53561 42517 53573 42520
rect 53607 42517 53619 42551
rect 55186 42548 55214 42588
rect 65794 42548 65800 42560
rect 55186 42520 65800 42548
rect 53561 42511 53619 42517
rect 65794 42508 65800 42520
rect 65852 42508 65858 42560
rect 552 42458 66424 42480
rect 552 42406 1998 42458
rect 2050 42406 2062 42458
rect 2114 42406 2126 42458
rect 2178 42406 2190 42458
rect 2242 42406 2254 42458
rect 2306 42406 50998 42458
rect 51050 42406 51062 42458
rect 51114 42406 51126 42458
rect 51178 42406 51190 42458
rect 51242 42406 51254 42458
rect 51306 42406 66424 42458
rect 552 42384 66424 42406
rect 10137 42347 10195 42353
rect 10137 42313 10149 42347
rect 10183 42344 10195 42347
rect 10410 42344 10416 42356
rect 10183 42316 10416 42344
rect 10183 42313 10195 42316
rect 10137 42307 10195 42313
rect 10410 42304 10416 42316
rect 10468 42344 10474 42356
rect 10468 42316 11652 42344
rect 10468 42304 10474 42316
rect 10229 42279 10287 42285
rect 10229 42245 10241 42279
rect 10275 42245 10287 42279
rect 10229 42239 10287 42245
rect 8665 42211 8723 42217
rect 8665 42177 8677 42211
rect 8711 42208 8723 42211
rect 10244 42208 10272 42239
rect 8711 42180 10272 42208
rect 8711 42177 8723 42180
rect 8665 42171 8723 42177
rect 10594 42168 10600 42220
rect 10652 42168 10658 42220
rect 10873 42211 10931 42217
rect 10873 42177 10885 42211
rect 10919 42208 10931 42211
rect 10962 42208 10968 42220
rect 10919 42180 10968 42208
rect 10919 42177 10931 42180
rect 10873 42171 10931 42177
rect 10962 42168 10968 42180
rect 11020 42168 11026 42220
rect 11624 42217 11652 42316
rect 13538 42304 13544 42356
rect 13596 42344 13602 42356
rect 15194 42344 15200 42356
rect 13596 42316 15200 42344
rect 13596 42304 13602 42316
rect 15194 42304 15200 42316
rect 15252 42304 15258 42356
rect 16022 42304 16028 42356
rect 16080 42344 16086 42356
rect 16482 42344 16488 42356
rect 16080 42316 16488 42344
rect 16080 42304 16086 42316
rect 16482 42304 16488 42316
rect 16540 42304 16546 42356
rect 16758 42304 16764 42356
rect 16816 42304 16822 42356
rect 20533 42347 20591 42353
rect 20533 42313 20545 42347
rect 20579 42344 20591 42347
rect 20714 42344 20720 42356
rect 20579 42316 20720 42344
rect 20579 42313 20591 42316
rect 20533 42307 20591 42313
rect 20714 42304 20720 42316
rect 20772 42304 20778 42356
rect 20806 42304 20812 42356
rect 20864 42344 20870 42356
rect 22094 42344 22100 42356
rect 20864 42316 22100 42344
rect 20864 42304 20870 42316
rect 22094 42304 22100 42316
rect 22152 42344 22158 42356
rect 22646 42344 22652 42356
rect 22152 42316 22652 42344
rect 22152 42304 22158 42316
rect 22646 42304 22652 42316
rect 22704 42344 22710 42356
rect 22704 42316 23980 42344
rect 22704 42304 22710 42316
rect 19613 42279 19671 42285
rect 19613 42276 19625 42279
rect 19076 42248 19625 42276
rect 11609 42211 11667 42217
rect 11609 42177 11621 42211
rect 11655 42177 11667 42211
rect 11609 42171 11667 42177
rect 14182 42168 14188 42220
rect 14240 42208 14246 42220
rect 14734 42208 14740 42220
rect 14240 42180 14740 42208
rect 14240 42168 14246 42180
rect 14734 42168 14740 42180
rect 14792 42168 14798 42220
rect 16666 42168 16672 42220
rect 16724 42208 16730 42220
rect 17405 42211 17463 42217
rect 17405 42208 17417 42211
rect 16724 42180 17417 42208
rect 16724 42168 16730 42180
rect 17405 42177 17417 42180
rect 17451 42208 17463 42211
rect 17862 42208 17868 42220
rect 17451 42180 17868 42208
rect 17451 42177 17463 42180
rect 17405 42171 17463 42177
rect 17862 42168 17868 42180
rect 17920 42168 17926 42220
rect 18046 42168 18052 42220
rect 18104 42168 18110 42220
rect 18233 42211 18291 42217
rect 18233 42177 18245 42211
rect 18279 42208 18291 42211
rect 18414 42208 18420 42220
rect 18279 42180 18420 42208
rect 18279 42177 18291 42180
rect 18233 42171 18291 42177
rect 18414 42168 18420 42180
rect 18472 42168 18478 42220
rect 7926 42100 7932 42152
rect 7984 42140 7990 42152
rect 8389 42143 8447 42149
rect 8389 42140 8401 42143
rect 7984 42112 8401 42140
rect 7984 42100 7990 42112
rect 8389 42109 8401 42112
rect 8435 42109 8447 42143
rect 8389 42103 8447 42109
rect 9766 42100 9772 42152
rect 9824 42140 9830 42152
rect 10612 42140 10640 42168
rect 9824 42112 10640 42140
rect 9824 42100 9830 42112
rect 17126 42100 17132 42152
rect 17184 42100 17190 42152
rect 18432 42140 18460 42168
rect 19076 42149 19104 42248
rect 19613 42245 19625 42248
rect 19659 42276 19671 42279
rect 23106 42276 23112 42288
rect 19659 42248 23112 42276
rect 19659 42245 19671 42248
rect 19613 42239 19671 42245
rect 23106 42236 23112 42248
rect 23164 42236 23170 42288
rect 23198 42236 23204 42288
rect 23256 42276 23262 42288
rect 23845 42279 23903 42285
rect 23845 42276 23857 42279
rect 23256 42248 23857 42276
rect 23256 42236 23262 42248
rect 23845 42245 23857 42248
rect 23891 42245 23903 42279
rect 23845 42239 23903 42245
rect 19150 42168 19156 42220
rect 19208 42168 19214 42220
rect 19242 42168 19248 42220
rect 19300 42168 19306 42220
rect 21818 42168 21824 42220
rect 21876 42208 21882 42220
rect 22554 42208 22560 42220
rect 21876 42180 22560 42208
rect 21876 42168 21882 42180
rect 22554 42168 22560 42180
rect 22612 42168 22618 42220
rect 23014 42168 23020 42220
rect 23072 42168 23078 42220
rect 23952 42208 23980 42316
rect 24578 42304 24584 42356
rect 24636 42344 24642 42356
rect 24673 42347 24731 42353
rect 24673 42344 24685 42347
rect 24636 42316 24685 42344
rect 24636 42304 24642 42316
rect 24673 42313 24685 42316
rect 24719 42313 24731 42347
rect 24673 42307 24731 42313
rect 25130 42304 25136 42356
rect 25188 42344 25194 42356
rect 25188 42316 26188 42344
rect 25188 42304 25194 42316
rect 24762 42236 24768 42288
rect 24820 42276 24826 42288
rect 25685 42279 25743 42285
rect 25685 42276 25697 42279
rect 24820 42248 25697 42276
rect 24820 42236 24826 42248
rect 25685 42245 25697 42248
rect 25731 42245 25743 42279
rect 25685 42239 25743 42245
rect 24397 42211 24455 42217
rect 24397 42208 24409 42211
rect 23952 42180 24409 42208
rect 24397 42177 24409 42180
rect 24443 42177 24455 42211
rect 24397 42171 24455 42177
rect 25038 42168 25044 42220
rect 25096 42208 25102 42220
rect 25133 42211 25191 42217
rect 25133 42208 25145 42211
rect 25096 42180 25145 42208
rect 25096 42168 25102 42180
rect 25133 42177 25145 42180
rect 25179 42177 25191 42211
rect 25133 42171 25191 42177
rect 25317 42211 25375 42217
rect 25317 42177 25329 42211
rect 25363 42208 25375 42211
rect 25958 42208 25964 42220
rect 25363 42180 25964 42208
rect 25363 42177 25375 42180
rect 25317 42171 25375 42177
rect 25958 42168 25964 42180
rect 26016 42168 26022 42220
rect 26160 42217 26188 42316
rect 26804 42316 28212 42344
rect 26145 42211 26203 42217
rect 26145 42177 26157 42211
rect 26191 42177 26203 42211
rect 26145 42171 26203 42177
rect 26234 42168 26240 42220
rect 26292 42168 26298 42220
rect 19061 42143 19119 42149
rect 18432 42112 19012 42140
rect 10597 42075 10655 42081
rect 10597 42041 10609 42075
rect 10643 42072 10655 42075
rect 11057 42075 11115 42081
rect 11057 42072 11069 42075
rect 10643 42044 11069 42072
rect 10643 42041 10655 42044
rect 10597 42035 10655 42041
rect 11057 42041 11069 42044
rect 11103 42041 11115 42075
rect 11057 42035 11115 42041
rect 15010 42032 15016 42084
rect 15068 42032 15074 42084
rect 16298 42072 16304 42084
rect 16238 42044 16304 42072
rect 16298 42032 16304 42044
rect 16356 42072 16362 42084
rect 16942 42072 16948 42084
rect 16356 42044 16948 42072
rect 16356 42032 16362 42044
rect 16942 42032 16948 42044
rect 17000 42032 17006 42084
rect 17221 42075 17279 42081
rect 17221 42041 17233 42075
rect 17267 42072 17279 42075
rect 18984 42072 19012 42112
rect 19061 42109 19073 42143
rect 19107 42109 19119 42143
rect 19260 42140 19288 42168
rect 19061 42103 19119 42109
rect 19168 42112 19288 42140
rect 19168 42072 19196 42112
rect 22922 42100 22928 42152
rect 22980 42140 22986 42152
rect 23293 42143 23351 42149
rect 23293 42140 23305 42143
rect 22980 42112 23305 42140
rect 22980 42100 22986 42112
rect 23293 42109 23305 42112
rect 23339 42109 23351 42143
rect 23293 42103 23351 42109
rect 24210 42100 24216 42152
rect 24268 42140 24274 42152
rect 24578 42140 24584 42152
rect 24268 42112 24584 42140
rect 24268 42100 24274 42112
rect 24578 42100 24584 42112
rect 24636 42100 24642 42152
rect 26804 42140 26832 42316
rect 26878 42168 26884 42220
rect 26936 42168 26942 42220
rect 27157 42211 27215 42217
rect 27157 42177 27169 42211
rect 27203 42208 27215 42211
rect 27614 42208 27620 42220
rect 27203 42180 27620 42208
rect 27203 42177 27215 42180
rect 27157 42171 27215 42177
rect 27614 42168 27620 42180
rect 27672 42168 27678 42220
rect 28184 42208 28212 42316
rect 28626 42304 28632 42356
rect 28684 42304 28690 42356
rect 28994 42304 29000 42356
rect 29052 42304 29058 42356
rect 33594 42304 33600 42356
rect 33652 42344 33658 42356
rect 34149 42347 34207 42353
rect 34149 42344 34161 42347
rect 33652 42316 34161 42344
rect 33652 42304 33658 42316
rect 34149 42313 34161 42316
rect 34195 42313 34207 42347
rect 34149 42307 34207 42313
rect 35066 42304 35072 42356
rect 35124 42304 35130 42356
rect 35158 42304 35164 42356
rect 35216 42344 35222 42356
rect 35253 42347 35311 42353
rect 35253 42344 35265 42347
rect 35216 42316 35265 42344
rect 35216 42304 35222 42316
rect 35253 42313 35265 42316
rect 35299 42313 35311 42347
rect 35253 42307 35311 42313
rect 36814 42304 36820 42356
rect 36872 42344 36878 42356
rect 37001 42347 37059 42353
rect 37001 42344 37013 42347
rect 36872 42316 37013 42344
rect 36872 42304 36878 42316
rect 37001 42313 37013 42316
rect 37047 42313 37059 42347
rect 37001 42307 37059 42313
rect 37292 42316 38516 42344
rect 28534 42236 28540 42288
rect 28592 42276 28598 42288
rect 30469 42279 30527 42285
rect 30469 42276 30481 42279
rect 28592 42248 30481 42276
rect 28592 42236 28598 42248
rect 30469 42245 30481 42248
rect 30515 42245 30527 42279
rect 30469 42239 30527 42245
rect 30834 42236 30840 42288
rect 30892 42276 30898 42288
rect 30892 42248 33824 42276
rect 30892 42236 30898 42248
rect 32306 42208 32312 42220
rect 28184 42180 32312 42208
rect 32306 42168 32312 42180
rect 32364 42168 32370 42220
rect 33134 42168 33140 42220
rect 33192 42208 33198 42220
rect 33410 42208 33416 42220
rect 33192 42180 33416 42208
rect 33192 42168 33198 42180
rect 33410 42168 33416 42180
rect 33468 42168 33474 42220
rect 26160 42112 26832 42140
rect 17267 42044 18736 42072
rect 18984 42044 19196 42072
rect 17267 42041 17279 42044
rect 17221 42035 17279 42041
rect 10686 41964 10692 42016
rect 10744 41964 10750 42016
rect 17589 42007 17647 42013
rect 17589 41973 17601 42007
rect 17635 42004 17647 42007
rect 17678 42004 17684 42016
rect 17635 41976 17684 42004
rect 17635 41973 17647 41976
rect 17589 41967 17647 41973
rect 17678 41964 17684 41976
rect 17736 41964 17742 42016
rect 17954 41964 17960 42016
rect 18012 41964 18018 42016
rect 18708 42013 18736 42044
rect 20530 42032 20536 42084
rect 20588 42072 20594 42084
rect 21821 42075 21879 42081
rect 21821 42072 21833 42075
rect 20588 42044 21833 42072
rect 20588 42032 20594 42044
rect 21821 42041 21833 42044
rect 21867 42072 21879 42075
rect 25774 42072 25780 42084
rect 21867 42044 25780 42072
rect 21867 42041 21879 42044
rect 21821 42035 21879 42041
rect 25774 42032 25780 42044
rect 25832 42032 25838 42084
rect 26053 42075 26111 42081
rect 26053 42041 26065 42075
rect 26099 42072 26111 42075
rect 26160 42072 26188 42112
rect 28258 42100 28264 42152
rect 28316 42100 28322 42152
rect 28626 42100 28632 42152
rect 28684 42140 28690 42152
rect 29549 42143 29607 42149
rect 29549 42140 29561 42143
rect 28684 42112 29561 42140
rect 28684 42100 28690 42112
rect 29549 42109 29561 42112
rect 29595 42109 29607 42143
rect 29549 42103 29607 42109
rect 30190 42100 30196 42152
rect 30248 42140 30254 42152
rect 32125 42143 32183 42149
rect 30248 42112 31754 42140
rect 30248 42100 30254 42112
rect 30650 42072 30656 42084
rect 26099 42044 26188 42072
rect 28460 42044 30656 42072
rect 26099 42041 26111 42044
rect 26053 42035 26111 42041
rect 18693 42007 18751 42013
rect 18693 41973 18705 42007
rect 18739 41973 18751 42007
rect 18693 41967 18751 41973
rect 22370 41964 22376 42016
rect 22428 41964 22434 42016
rect 23198 41964 23204 42016
rect 23256 41964 23262 42016
rect 23661 42007 23719 42013
rect 23661 41973 23673 42007
rect 23707 42004 23719 42007
rect 24118 42004 24124 42016
rect 23707 41976 24124 42004
rect 23707 41973 23719 41976
rect 23661 41967 23719 41973
rect 24118 41964 24124 41976
rect 24176 41964 24182 42016
rect 24210 41964 24216 42016
rect 24268 42004 24274 42016
rect 24305 42007 24363 42013
rect 24305 42004 24317 42007
rect 24268 41976 24317 42004
rect 24268 41964 24274 41976
rect 24305 41973 24317 41976
rect 24351 41973 24363 42007
rect 24305 41967 24363 41973
rect 25041 42007 25099 42013
rect 25041 41973 25053 42007
rect 25087 42004 25099 42007
rect 25406 42004 25412 42016
rect 25087 41976 25412 42004
rect 25087 41973 25099 41976
rect 25041 41967 25099 41973
rect 25406 41964 25412 41976
rect 25464 41964 25470 42016
rect 25593 42007 25651 42013
rect 25593 41973 25605 42007
rect 25639 42004 25651 42007
rect 25866 42004 25872 42016
rect 25639 41976 25872 42004
rect 25639 41973 25651 41976
rect 25593 41967 25651 41973
rect 25866 41964 25872 41976
rect 25924 42004 25930 42016
rect 28460 42004 28488 42044
rect 30650 42032 30656 42044
rect 30708 42032 30714 42084
rect 30742 42032 30748 42084
rect 30800 42032 30806 42084
rect 31726 42072 31754 42112
rect 32125 42109 32137 42143
rect 32171 42140 32183 42143
rect 33686 42140 33692 42152
rect 32171 42112 33692 42140
rect 32171 42109 32183 42112
rect 32125 42103 32183 42109
rect 33686 42100 33692 42112
rect 33744 42100 33750 42152
rect 33796 42149 33824 42248
rect 34790 42236 34796 42288
rect 34848 42276 34854 42288
rect 37292 42276 37320 42316
rect 34848 42248 37320 42276
rect 38488 42276 38516 42316
rect 38930 42304 38936 42356
rect 38988 42344 38994 42356
rect 39298 42344 39304 42356
rect 38988 42316 39304 42344
rect 38988 42304 38994 42316
rect 39298 42304 39304 42316
rect 39356 42304 39362 42356
rect 42058 42304 42064 42356
rect 42116 42304 42122 42356
rect 51626 42344 51632 42356
rect 43732 42316 51632 42344
rect 38488 42248 40724 42276
rect 34848 42236 34854 42248
rect 34606 42168 34612 42220
rect 34664 42168 34670 42220
rect 34701 42211 34759 42217
rect 34701 42177 34713 42211
rect 34747 42177 34759 42211
rect 34701 42171 34759 42177
rect 33781 42143 33839 42149
rect 33781 42109 33793 42143
rect 33827 42109 33839 42143
rect 33781 42103 33839 42109
rect 33965 42143 34023 42149
rect 33965 42109 33977 42143
rect 34011 42140 34023 42143
rect 34011 42112 34376 42140
rect 34011 42109 34023 42112
rect 33965 42103 34023 42109
rect 31846 42072 31852 42084
rect 31726 42044 31852 42072
rect 31846 42032 31852 42044
rect 31904 42032 31910 42084
rect 32398 42072 32404 42084
rect 31956 42044 32404 42072
rect 25924 41976 28488 42004
rect 30285 42007 30343 42013
rect 25924 41964 25930 41976
rect 30285 41973 30297 42007
rect 30331 42004 30343 42007
rect 30374 42004 30380 42016
rect 30331 41976 30380 42004
rect 30331 41973 30343 41976
rect 30285 41967 30343 41973
rect 30374 41964 30380 41976
rect 30432 41964 30438 42016
rect 30466 41964 30472 42016
rect 30524 42004 30530 42016
rect 31956 42004 31984 42044
rect 32398 42032 32404 42044
rect 32456 42032 32462 42084
rect 32677 42075 32735 42081
rect 32677 42041 32689 42075
rect 32723 42072 32735 42075
rect 32723 42044 32996 42072
rect 32723 42041 32735 42044
rect 32677 42035 32735 42041
rect 30524 41976 31984 42004
rect 30524 41964 30530 41976
rect 32214 41964 32220 42016
rect 32272 42004 32278 42016
rect 32769 42007 32827 42013
rect 32769 42004 32781 42007
rect 32272 41976 32781 42004
rect 32272 41964 32278 41976
rect 32769 41973 32781 41976
rect 32815 41973 32827 42007
rect 32968 42004 32996 42044
rect 33410 42032 33416 42084
rect 33468 42072 33474 42084
rect 34238 42072 34244 42084
rect 33468 42044 34244 42072
rect 33468 42032 33474 42044
rect 34238 42032 34244 42044
rect 34296 42032 34302 42084
rect 34348 42072 34376 42112
rect 34422 42100 34428 42152
rect 34480 42140 34486 42152
rect 34716 42140 34744 42171
rect 35710 42168 35716 42220
rect 35768 42168 35774 42220
rect 35802 42168 35808 42220
rect 35860 42168 35866 42220
rect 37461 42211 37519 42217
rect 37461 42177 37473 42211
rect 37507 42208 37519 42211
rect 37826 42208 37832 42220
rect 37507 42180 37832 42208
rect 37507 42177 37519 42180
rect 37461 42171 37519 42177
rect 37826 42168 37832 42180
rect 37884 42168 37890 42220
rect 34480 42112 34744 42140
rect 35621 42143 35679 42149
rect 34480 42100 34486 42112
rect 35621 42109 35633 42143
rect 35667 42140 35679 42143
rect 35894 42140 35900 42152
rect 35667 42112 35900 42140
rect 35667 42109 35679 42112
rect 35621 42103 35679 42109
rect 35894 42100 35900 42112
rect 35952 42100 35958 42152
rect 36081 42143 36139 42149
rect 36081 42109 36093 42143
rect 36127 42140 36139 42143
rect 36262 42140 36268 42152
rect 36127 42112 36268 42140
rect 36127 42109 36139 42112
rect 36081 42103 36139 42109
rect 36262 42100 36268 42112
rect 36320 42140 36326 42152
rect 37185 42143 37243 42149
rect 37185 42140 37197 42143
rect 36320 42112 37197 42140
rect 36320 42100 36326 42112
rect 37185 42109 37197 42112
rect 37231 42109 37243 42143
rect 37185 42103 37243 42109
rect 39945 42143 40003 42149
rect 39945 42109 39957 42143
rect 39991 42140 40003 42143
rect 40034 42140 40040 42152
rect 39991 42112 40040 42140
rect 39991 42109 40003 42112
rect 39945 42103 40003 42109
rect 40034 42100 40040 42112
rect 40092 42100 40098 42152
rect 40696 42140 40724 42248
rect 40862 42236 40868 42288
rect 40920 42276 40926 42288
rect 40920 42248 43024 42276
rect 40920 42236 40926 42248
rect 40773 42211 40831 42217
rect 40773 42177 40785 42211
rect 40819 42208 40831 42211
rect 41598 42208 41604 42220
rect 40819 42180 41604 42208
rect 40819 42177 40831 42180
rect 40773 42171 40831 42177
rect 41598 42168 41604 42180
rect 41656 42208 41662 42220
rect 42426 42208 42432 42220
rect 41656 42180 42432 42208
rect 41656 42168 41662 42180
rect 42426 42168 42432 42180
rect 42484 42168 42490 42220
rect 42610 42168 42616 42220
rect 42668 42168 42674 42220
rect 40696 42112 41184 42140
rect 34974 42072 34980 42084
rect 34348 42044 34980 42072
rect 34974 42032 34980 42044
rect 35032 42032 35038 42084
rect 38746 42072 38752 42084
rect 38686 42044 38752 42072
rect 38746 42032 38752 42044
rect 38804 42072 38810 42084
rect 39390 42072 39396 42084
rect 38804 42044 39396 42072
rect 38804 42032 38810 42044
rect 39390 42032 39396 42044
rect 39448 42032 39454 42084
rect 40589 42075 40647 42081
rect 40589 42041 40601 42075
rect 40635 42072 40647 42075
rect 41049 42075 41107 42081
rect 41049 42072 41061 42075
rect 40635 42044 41061 42072
rect 40635 42041 40647 42044
rect 40589 42035 40647 42041
rect 41049 42041 41061 42044
rect 41095 42041 41107 42075
rect 41156 42072 41184 42112
rect 41690 42100 41696 42152
rect 41748 42100 41754 42152
rect 42521 42143 42579 42149
rect 42521 42109 42533 42143
rect 42567 42140 42579 42143
rect 42702 42140 42708 42152
rect 42567 42112 42708 42140
rect 42567 42109 42579 42112
rect 42521 42103 42579 42109
rect 42702 42100 42708 42112
rect 42760 42100 42766 42152
rect 42996 42149 43024 42248
rect 43346 42236 43352 42288
rect 43404 42276 43410 42288
rect 43441 42279 43499 42285
rect 43441 42276 43453 42279
rect 43404 42248 43453 42276
rect 43404 42236 43410 42248
rect 43441 42245 43453 42248
rect 43487 42245 43499 42279
rect 43441 42239 43499 42245
rect 42981 42143 43039 42149
rect 42981 42109 42993 42143
rect 43027 42140 43039 42143
rect 43732 42140 43760 42316
rect 51626 42304 51632 42316
rect 51684 42304 51690 42356
rect 51718 42304 51724 42356
rect 51776 42344 51782 42356
rect 51776 42316 53972 42344
rect 51776 42304 51782 42316
rect 43898 42236 43904 42288
rect 43956 42276 43962 42288
rect 43956 42248 44956 42276
rect 43956 42236 43962 42248
rect 43990 42168 43996 42220
rect 44048 42168 44054 42220
rect 44928 42217 44956 42248
rect 44913 42211 44971 42217
rect 44913 42177 44925 42211
rect 44959 42177 44971 42211
rect 44913 42171 44971 42177
rect 45005 42211 45063 42217
rect 45005 42177 45017 42211
rect 45051 42177 45063 42211
rect 45005 42171 45063 42177
rect 43027 42112 43760 42140
rect 43809 42143 43867 42149
rect 43027 42109 43039 42112
rect 42981 42103 43039 42109
rect 43809 42109 43821 42143
rect 43855 42140 43867 42143
rect 44082 42140 44088 42152
rect 43855 42112 44088 42140
rect 43855 42109 43867 42112
rect 43809 42103 43867 42109
rect 44082 42100 44088 42112
rect 44140 42100 44146 42152
rect 44174 42100 44180 42152
rect 44232 42140 44238 42152
rect 45020 42140 45048 42171
rect 45462 42168 45468 42220
rect 45520 42208 45526 42220
rect 46934 42208 46940 42220
rect 45520 42180 46940 42208
rect 45520 42168 45526 42180
rect 46934 42168 46940 42180
rect 46992 42168 46998 42220
rect 47305 42211 47363 42217
rect 47305 42177 47317 42211
rect 47351 42208 47363 42211
rect 47394 42208 47400 42220
rect 47351 42180 47400 42208
rect 47351 42177 47363 42180
rect 47305 42171 47363 42177
rect 47394 42168 47400 42180
rect 47452 42168 47458 42220
rect 47670 42168 47676 42220
rect 47728 42168 47734 42220
rect 48682 42168 48688 42220
rect 48740 42208 48746 42220
rect 49050 42208 49056 42220
rect 48740 42180 49056 42208
rect 48740 42168 48746 42180
rect 49050 42168 49056 42180
rect 49108 42208 49114 42220
rect 49421 42211 49479 42217
rect 49421 42208 49433 42211
rect 49108 42180 49433 42208
rect 49108 42168 49114 42180
rect 49421 42177 49433 42180
rect 49467 42177 49479 42211
rect 49421 42171 49479 42177
rect 51350 42168 51356 42220
rect 51408 42208 51414 42220
rect 52641 42211 52699 42217
rect 52641 42208 52653 42211
rect 51408 42180 52653 42208
rect 51408 42168 51414 42180
rect 52641 42177 52653 42180
rect 52687 42177 52699 42211
rect 52641 42171 52699 42177
rect 53377 42211 53435 42217
rect 53377 42177 53389 42211
rect 53423 42208 53435 42211
rect 53423 42180 53880 42208
rect 53423 42177 53435 42180
rect 53377 42171 53435 42177
rect 44232 42112 45048 42140
rect 44232 42100 44238 42112
rect 53098 42100 53104 42152
rect 53156 42100 53162 42152
rect 41156 42044 41414 42072
rect 41049 42035 41107 42041
rect 33137 42007 33195 42013
rect 33137 42004 33149 42007
rect 32968 41976 33149 42004
rect 32769 41967 32827 41973
rect 33137 41973 33149 41976
rect 33183 41973 33195 42007
rect 33137 41967 33195 41973
rect 33226 41964 33232 42016
rect 33284 41964 33290 42016
rect 33318 41964 33324 42016
rect 33376 42004 33382 42016
rect 34517 42007 34575 42013
rect 34517 42004 34529 42007
rect 33376 41976 34529 42004
rect 33376 41964 33382 41976
rect 34517 41973 34529 41976
rect 34563 41973 34575 42007
rect 34517 41967 34575 41973
rect 39298 41964 39304 42016
rect 39356 41964 39362 42016
rect 39850 41964 39856 42016
rect 39908 42004 39914 42016
rect 40221 42007 40279 42013
rect 40221 42004 40233 42007
rect 39908 41976 40233 42004
rect 39908 41964 39914 41976
rect 40221 41973 40233 41976
rect 40267 41973 40279 42007
rect 40221 41967 40279 41973
rect 40310 41964 40316 42016
rect 40368 42004 40374 42016
rect 40681 42007 40739 42013
rect 40681 42004 40693 42007
rect 40368 41976 40693 42004
rect 40368 41964 40374 41976
rect 40681 41973 40693 41976
rect 40727 41973 40739 42007
rect 41386 42004 41414 42044
rect 41874 42032 41880 42084
rect 41932 42072 41938 42084
rect 42429 42075 42487 42081
rect 42429 42072 42441 42075
rect 41932 42044 42441 42072
rect 41932 42032 41938 42044
rect 42429 42041 42441 42044
rect 42475 42041 42487 42075
rect 42429 42035 42487 42041
rect 43349 42075 43407 42081
rect 43349 42041 43361 42075
rect 43395 42072 43407 42075
rect 43438 42072 43444 42084
rect 43395 42044 43444 42072
rect 43395 42041 43407 42044
rect 43349 42035 43407 42041
rect 43438 42032 43444 42044
rect 43496 42032 43502 42084
rect 43622 42032 43628 42084
rect 43680 42072 43686 42084
rect 43901 42075 43959 42081
rect 43901 42072 43913 42075
rect 43680 42044 43913 42072
rect 43680 42032 43686 42044
rect 43901 42041 43913 42044
rect 43947 42041 43959 42075
rect 45281 42075 45339 42081
rect 45281 42072 45293 42075
rect 43901 42035 43959 42041
rect 44836 42044 45293 42072
rect 44836 42016 44864 42044
rect 45281 42041 45293 42044
rect 45327 42041 45339 42075
rect 45281 42035 45339 42041
rect 46014 42032 46020 42084
rect 46072 42032 46078 42084
rect 47026 42032 47032 42084
rect 47084 42032 47090 42084
rect 48130 42032 48136 42084
rect 48188 42032 48194 42084
rect 50614 42032 50620 42084
rect 50672 42032 50678 42084
rect 51810 42032 51816 42084
rect 51868 42032 51874 42084
rect 52365 42075 52423 42081
rect 52365 42041 52377 42075
rect 52411 42072 52423 42075
rect 53852 42072 53880 42180
rect 53944 42149 53972 42316
rect 54202 42168 54208 42220
rect 54260 42168 54266 42220
rect 53929 42143 53987 42149
rect 53929 42109 53941 42143
rect 53975 42109 53987 42143
rect 53929 42103 53987 42109
rect 54018 42100 54024 42152
rect 54076 42140 54082 42152
rect 55033 42143 55091 42149
rect 55033 42140 55045 42143
rect 54076 42112 55045 42140
rect 54076 42100 54082 42112
rect 55033 42109 55045 42112
rect 55079 42140 55091 42143
rect 63034 42140 63040 42152
rect 55079 42112 63040 42140
rect 55079 42109 55091 42112
rect 55033 42103 55091 42109
rect 63034 42100 63040 42112
rect 63092 42100 63098 42152
rect 54478 42072 54484 42084
rect 52411 42044 53604 42072
rect 53852 42044 54484 42072
rect 52411 42041 52423 42044
rect 52365 42035 52423 42041
rect 43070 42004 43076 42016
rect 41386 41976 43076 42004
rect 40681 41967 40739 41973
rect 43070 41964 43076 41976
rect 43128 41964 43134 42016
rect 44450 41964 44456 42016
rect 44508 41964 44514 42016
rect 44818 41964 44824 42016
rect 44876 41964 44882 42016
rect 45554 41964 45560 42016
rect 45612 42004 45618 42016
rect 46842 42004 46848 42016
rect 45612 41976 46848 42004
rect 45612 41964 45618 41976
rect 46842 41964 46848 41976
rect 46900 41964 46906 42016
rect 46934 41964 46940 42016
rect 46992 42004 46998 42016
rect 52270 42004 52276 42016
rect 46992 41976 52276 42004
rect 46992 41964 46998 41976
rect 52270 41964 52276 41976
rect 52328 41964 52334 42016
rect 52454 41964 52460 42016
rect 52512 42004 52518 42016
rect 52733 42007 52791 42013
rect 52733 42004 52745 42007
rect 52512 41976 52745 42004
rect 52512 41964 52518 41976
rect 52733 41973 52745 41976
rect 52779 41973 52791 42007
rect 52733 41967 52791 41973
rect 53190 41964 53196 42016
rect 53248 41964 53254 42016
rect 53576 42013 53604 42044
rect 54478 42032 54484 42044
rect 54536 42032 54542 42084
rect 53561 42007 53619 42013
rect 53561 41973 53573 42007
rect 53607 41973 53619 42007
rect 53561 41967 53619 41973
rect 54018 41964 54024 42016
rect 54076 41964 54082 42016
rect 54846 41964 54852 42016
rect 54904 41964 54910 42016
rect 552 41914 66424 41936
rect 552 41862 2918 41914
rect 2970 41862 2982 41914
rect 3034 41862 3046 41914
rect 3098 41862 3110 41914
rect 3162 41862 3174 41914
rect 3226 41862 51918 41914
rect 51970 41862 51982 41914
rect 52034 41862 52046 41914
rect 52098 41862 52110 41914
rect 52162 41862 52174 41914
rect 52226 41862 66424 41914
rect 552 41840 66424 41862
rect 10410 41760 10416 41812
rect 10468 41760 10474 41812
rect 15010 41760 15016 41812
rect 15068 41800 15074 41812
rect 15197 41803 15255 41809
rect 15197 41800 15209 41803
rect 15068 41772 15209 41800
rect 15068 41760 15074 41772
rect 15197 41769 15209 41772
rect 15243 41769 15255 41803
rect 15197 41763 15255 41769
rect 15562 41760 15568 41812
rect 15620 41760 15626 41812
rect 15657 41803 15715 41809
rect 15657 41769 15669 41803
rect 15703 41800 15715 41803
rect 16393 41803 16451 41809
rect 16393 41800 16405 41803
rect 15703 41772 16405 41800
rect 15703 41769 15715 41772
rect 15657 41763 15715 41769
rect 16393 41769 16405 41772
rect 16439 41769 16451 41803
rect 16393 41763 16451 41769
rect 16574 41760 16580 41812
rect 16632 41800 16638 41812
rect 17221 41803 17279 41809
rect 17221 41800 17233 41803
rect 16632 41772 17233 41800
rect 16632 41760 16638 41772
rect 17221 41769 17233 41772
rect 17267 41769 17279 41803
rect 17221 41763 17279 41769
rect 17586 41760 17592 41812
rect 17644 41760 17650 41812
rect 17678 41760 17684 41812
rect 17736 41760 17742 41812
rect 20714 41760 20720 41812
rect 20772 41760 20778 41812
rect 23474 41800 23480 41812
rect 21284 41772 23480 41800
rect 9766 41732 9772 41744
rect 9430 41704 9772 41732
rect 9766 41692 9772 41704
rect 9824 41692 9830 41744
rect 15378 41692 15384 41744
rect 15436 41732 15442 41744
rect 16853 41735 16911 41741
rect 16853 41732 16865 41735
rect 15436 41704 16865 41732
rect 15436 41692 15442 41704
rect 16853 41701 16865 41704
rect 16899 41732 16911 41735
rect 17954 41732 17960 41744
rect 16899 41704 17960 41732
rect 16899 41701 16911 41704
rect 16853 41695 16911 41701
rect 17954 41692 17960 41704
rect 18012 41692 18018 41744
rect 20732 41732 20760 41760
rect 21284 41732 21312 41772
rect 23474 41760 23480 41772
rect 23532 41800 23538 41812
rect 23658 41800 23664 41812
rect 23532 41772 23664 41800
rect 23532 41760 23538 41772
rect 23658 41760 23664 41772
rect 23716 41760 23722 41812
rect 23842 41760 23848 41812
rect 23900 41800 23906 41812
rect 23900 41772 25728 41800
rect 23900 41760 23906 41772
rect 20732 41704 21312 41732
rect 10505 41667 10563 41673
rect 10505 41633 10517 41667
rect 10551 41664 10563 41667
rect 11422 41664 11428 41676
rect 10551 41636 11428 41664
rect 10551 41633 10563 41636
rect 10505 41627 10563 41633
rect 11422 41624 11428 41636
rect 11480 41624 11486 41676
rect 12713 41667 12771 41673
rect 12713 41633 12725 41667
rect 12759 41664 12771 41667
rect 13173 41667 13231 41673
rect 13173 41664 13185 41667
rect 12759 41636 13185 41664
rect 12759 41633 12771 41636
rect 12713 41627 12771 41633
rect 13173 41633 13185 41636
rect 13219 41633 13231 41667
rect 13173 41627 13231 41633
rect 14277 41667 14335 41673
rect 14277 41633 14289 41667
rect 14323 41633 14335 41667
rect 16666 41664 16672 41676
rect 14277 41627 14335 41633
rect 15856 41636 16672 41664
rect 7926 41556 7932 41608
rect 7984 41556 7990 41608
rect 8202 41556 8208 41608
rect 8260 41556 8266 41608
rect 10410 41556 10416 41608
rect 10468 41596 10474 41608
rect 10597 41599 10655 41605
rect 10597 41596 10609 41599
rect 10468 41568 10609 41596
rect 10468 41556 10474 41568
rect 10597 41565 10609 41568
rect 10643 41565 10655 41599
rect 10597 41559 10655 41565
rect 11330 41556 11336 41608
rect 11388 41596 11394 41608
rect 12161 41599 12219 41605
rect 12161 41596 12173 41599
rect 11388 41568 12173 41596
rect 11388 41556 11394 41568
rect 12161 41565 12173 41568
rect 12207 41565 12219 41599
rect 12161 41559 12219 41565
rect 12618 41556 12624 41608
rect 12676 41596 12682 41608
rect 12805 41599 12863 41605
rect 12805 41596 12817 41599
rect 12676 41568 12817 41596
rect 12676 41556 12682 41568
rect 12805 41565 12817 41568
rect 12851 41565 12863 41599
rect 12805 41559 12863 41565
rect 12894 41556 12900 41608
rect 12952 41556 12958 41608
rect 13814 41556 13820 41608
rect 13872 41556 13878 41608
rect 10962 41488 10968 41540
rect 11020 41528 11026 41540
rect 12912 41528 12940 41556
rect 13170 41528 13176 41540
rect 11020 41500 13176 41528
rect 11020 41488 11026 41500
rect 13170 41488 13176 41500
rect 13228 41488 13234 41540
rect 14292 41528 14320 41627
rect 15856 41605 15884 41636
rect 16666 41624 16672 41636
rect 16724 41624 16730 41676
rect 16758 41624 16764 41676
rect 16816 41624 16822 41676
rect 21284 41673 21312 41704
rect 22186 41692 22192 41744
rect 22244 41692 22250 41744
rect 23109 41735 23167 41741
rect 23109 41701 23121 41735
rect 23155 41732 23167 41735
rect 23382 41732 23388 41744
rect 23155 41704 23388 41732
rect 23155 41701 23167 41704
rect 23109 41695 23167 41701
rect 23382 41692 23388 41704
rect 23440 41692 23446 41744
rect 24210 41732 24216 41744
rect 23492 41704 24216 41732
rect 19521 41667 19579 41673
rect 19521 41633 19533 41667
rect 19567 41664 19579 41667
rect 20717 41667 20775 41673
rect 20717 41664 20729 41667
rect 19567 41636 20729 41664
rect 19567 41633 19579 41636
rect 19521 41627 19579 41633
rect 20717 41633 20729 41636
rect 20763 41633 20775 41667
rect 20717 41627 20775 41633
rect 21269 41667 21327 41673
rect 21269 41633 21281 41667
rect 21315 41633 21327 41667
rect 21269 41627 21327 41633
rect 15841 41599 15899 41605
rect 15841 41565 15853 41599
rect 15887 41565 15899 41599
rect 15841 41559 15899 41565
rect 16390 41556 16396 41608
rect 16448 41596 16454 41608
rect 16945 41599 17003 41605
rect 16945 41596 16957 41599
rect 16448 41568 16957 41596
rect 16448 41556 16454 41568
rect 16945 41565 16957 41568
rect 16991 41565 17003 41599
rect 16945 41559 17003 41565
rect 17862 41556 17868 41608
rect 17920 41556 17926 41608
rect 18322 41556 18328 41608
rect 18380 41596 18386 41608
rect 18601 41599 18659 41605
rect 18601 41596 18613 41599
rect 18380 41568 18613 41596
rect 18380 41556 18386 41568
rect 18601 41565 18613 41568
rect 18647 41565 18659 41599
rect 18601 41559 18659 41565
rect 18969 41599 19027 41605
rect 18969 41565 18981 41599
rect 19015 41565 19027 41599
rect 18969 41559 19027 41565
rect 20257 41599 20315 41605
rect 20257 41565 20269 41599
rect 20303 41596 20315 41599
rect 20622 41596 20628 41608
rect 20303 41568 20628 41596
rect 20303 41565 20315 41568
rect 20257 41559 20315 41565
rect 18874 41528 18880 41540
rect 14292 41500 18880 41528
rect 18874 41488 18880 41500
rect 18932 41488 18938 41540
rect 18984 41528 19012 41559
rect 20622 41556 20628 41568
rect 20680 41556 20686 41608
rect 20809 41599 20867 41605
rect 20809 41565 20821 41599
rect 20855 41565 20867 41599
rect 20809 41559 20867 41565
rect 20824 41528 20852 41559
rect 20990 41556 20996 41608
rect 21048 41556 21054 41608
rect 21542 41556 21548 41608
rect 21600 41556 21606 41608
rect 22830 41556 22836 41608
rect 22888 41596 22894 41608
rect 23017 41599 23075 41605
rect 23017 41596 23029 41599
rect 22888 41568 23029 41596
rect 22888 41556 22894 41568
rect 23017 41565 23029 41568
rect 23063 41596 23075 41599
rect 23492 41596 23520 41704
rect 24210 41692 24216 41704
rect 24268 41692 24274 41744
rect 24854 41692 24860 41744
rect 24912 41692 24918 41744
rect 25700 41741 25728 41772
rect 25774 41760 25780 41812
rect 25832 41800 25838 41812
rect 27062 41800 27068 41812
rect 25832 41772 27068 41800
rect 25832 41760 25838 41772
rect 27062 41760 27068 41772
rect 27120 41760 27126 41812
rect 27522 41760 27528 41812
rect 27580 41800 27586 41812
rect 27580 41772 28028 41800
rect 27580 41760 27586 41772
rect 25685 41735 25743 41741
rect 25685 41701 25697 41735
rect 25731 41701 25743 41735
rect 25685 41695 25743 41701
rect 23842 41624 23848 41676
rect 23900 41624 23906 41676
rect 25700 41664 25728 41695
rect 26694 41692 26700 41744
rect 26752 41692 26758 41744
rect 28000 41732 28028 41772
rect 28166 41760 28172 41812
rect 28224 41800 28230 41812
rect 28629 41803 28687 41809
rect 28629 41800 28641 41803
rect 28224 41772 28641 41800
rect 28224 41760 28230 41772
rect 28629 41769 28641 41772
rect 28675 41769 28687 41803
rect 28629 41763 28687 41769
rect 28736 41772 33548 41800
rect 28736 41732 28764 41772
rect 28000 41704 28764 41732
rect 28997 41735 29055 41741
rect 28997 41701 29009 41735
rect 29043 41732 29055 41735
rect 30834 41732 30840 41744
rect 29043 41704 30840 41732
rect 29043 41701 29055 41704
rect 28997 41695 29055 41701
rect 30834 41692 30840 41704
rect 30892 41692 30898 41744
rect 32214 41692 32220 41744
rect 32272 41692 32278 41744
rect 33520 41732 33548 41772
rect 33686 41760 33692 41812
rect 33744 41760 33750 41812
rect 37185 41803 37243 41809
rect 37185 41769 37197 41803
rect 37231 41800 37243 41803
rect 39298 41800 39304 41812
rect 37231 41772 39304 41800
rect 37231 41769 37243 41772
rect 37185 41763 37243 41769
rect 39298 41760 39304 41772
rect 39356 41760 39362 41812
rect 40218 41760 40224 41812
rect 40276 41760 40282 41812
rect 41325 41803 41383 41809
rect 41325 41769 41337 41803
rect 41371 41800 41383 41803
rect 41690 41800 41696 41812
rect 41371 41772 41696 41800
rect 41371 41769 41383 41772
rect 41325 41763 41383 41769
rect 41690 41760 41696 41772
rect 41748 41800 41754 41812
rect 42429 41803 42487 41809
rect 42429 41800 42441 41803
rect 41748 41772 42441 41800
rect 41748 41760 41754 41772
rect 42429 41769 42441 41772
rect 42475 41769 42487 41803
rect 42429 41763 42487 41769
rect 42518 41760 42524 41812
rect 42576 41800 42582 41812
rect 44729 41803 44787 41809
rect 42576 41772 44588 41800
rect 42576 41760 42582 41772
rect 36998 41732 37004 41744
rect 33520 41704 37004 41732
rect 36998 41692 37004 41704
rect 37056 41692 37062 41744
rect 37090 41692 37096 41744
rect 37148 41732 37154 41744
rect 37645 41735 37703 41741
rect 37645 41732 37657 41735
rect 37148 41704 37657 41732
rect 37148 41692 37154 41704
rect 37645 41701 37657 41704
rect 37691 41701 37703 41735
rect 37645 41695 37703 41701
rect 38562 41692 38568 41744
rect 38620 41732 38626 41744
rect 39393 41735 39451 41741
rect 39393 41732 39405 41735
rect 38620 41704 39405 41732
rect 38620 41692 38626 41704
rect 39393 41701 39405 41704
rect 39439 41701 39451 41735
rect 40236 41732 40264 41760
rect 39393 41695 39451 41701
rect 39592 41704 40264 41732
rect 43257 41735 43315 41741
rect 26234 41664 26240 41676
rect 25700 41636 26240 41664
rect 26234 41624 26240 41636
rect 26292 41664 26298 41676
rect 26421 41667 26479 41673
rect 26421 41664 26433 41667
rect 26292 41636 26433 41664
rect 26292 41624 26298 41636
rect 26421 41633 26433 41636
rect 26467 41633 26479 41667
rect 28534 41664 28540 41676
rect 27830 41650 28540 41664
rect 26421 41627 26479 41633
rect 27816 41636 28540 41650
rect 23063 41568 23520 41596
rect 23063 41565 23075 41568
rect 23017 41559 23075 41565
rect 23750 41556 23756 41608
rect 23808 41556 23814 41608
rect 24118 41556 24124 41608
rect 24176 41556 24182 41608
rect 25130 41556 25136 41608
rect 25188 41596 25194 41608
rect 25593 41599 25651 41605
rect 25593 41596 25605 41599
rect 25188 41568 25605 41596
rect 25188 41556 25194 41568
rect 25593 41565 25605 41568
rect 25639 41565 25651 41599
rect 27816 41596 27844 41636
rect 28534 41624 28540 41636
rect 28592 41624 28598 41676
rect 30098 41624 30104 41676
rect 30156 41664 30162 41676
rect 30193 41667 30251 41673
rect 30193 41664 30205 41667
rect 30156 41636 30205 41664
rect 30156 41624 30162 41636
rect 30193 41633 30205 41636
rect 30239 41633 30251 41667
rect 30193 41627 30251 41633
rect 33318 41624 33324 41676
rect 33376 41664 33382 41676
rect 34054 41664 34060 41676
rect 33376 41636 34060 41664
rect 33376 41624 33382 41636
rect 34054 41624 34060 41636
rect 34112 41624 34118 41676
rect 34974 41624 34980 41676
rect 35032 41664 35038 41676
rect 35069 41667 35127 41673
rect 35069 41664 35081 41667
rect 35032 41636 35081 41664
rect 35032 41624 35038 41636
rect 35069 41633 35081 41636
rect 35115 41633 35127 41667
rect 38378 41664 38384 41676
rect 35069 41627 35127 41633
rect 37016 41636 38384 41664
rect 25593 41559 25651 41565
rect 26252 41568 27844 41596
rect 28169 41599 28227 41605
rect 21266 41528 21272 41540
rect 18984 41500 20760 41528
rect 20824 41500 21272 41528
rect 9674 41420 9680 41472
rect 9732 41420 9738 41472
rect 10042 41420 10048 41472
rect 10100 41420 10106 41472
rect 10778 41420 10784 41472
rect 10836 41460 10842 41472
rect 11609 41463 11667 41469
rect 11609 41460 11621 41463
rect 10836 41432 11621 41460
rect 10836 41420 10842 41432
rect 11609 41429 11621 41432
rect 11655 41429 11667 41463
rect 11609 41423 11667 41429
rect 11882 41420 11888 41472
rect 11940 41460 11946 41472
rect 12345 41463 12403 41469
rect 12345 41460 12357 41463
rect 11940 41432 12357 41460
rect 11940 41420 11946 41432
rect 12345 41429 12357 41432
rect 12391 41429 12403 41463
rect 12345 41423 12403 41429
rect 14185 41463 14243 41469
rect 14185 41429 14197 41463
rect 14231 41460 14243 41463
rect 14642 41460 14648 41472
rect 14231 41432 14648 41460
rect 14231 41429 14243 41432
rect 14185 41423 14243 41429
rect 14642 41420 14648 41432
rect 14700 41420 14706 41472
rect 15378 41420 15384 41472
rect 15436 41460 15442 41472
rect 16390 41460 16396 41472
rect 15436 41432 16396 41460
rect 15436 41420 15442 41432
rect 16390 41420 16396 41432
rect 16448 41420 16454 41472
rect 18046 41420 18052 41472
rect 18104 41420 18110 41472
rect 19610 41420 19616 41472
rect 19668 41420 19674 41472
rect 20254 41420 20260 41472
rect 20312 41460 20318 41472
rect 20349 41463 20407 41469
rect 20349 41460 20361 41463
rect 20312 41432 20361 41460
rect 20312 41420 20318 41432
rect 20349 41429 20361 41432
rect 20395 41429 20407 41463
rect 20732 41460 20760 41500
rect 21266 41488 21272 41500
rect 21324 41488 21330 41540
rect 25866 41488 25872 41540
rect 25924 41528 25930 41540
rect 26252 41528 26280 41568
rect 28169 41565 28181 41599
rect 28215 41596 28227 41599
rect 28442 41596 28448 41608
rect 28215 41568 28448 41596
rect 28215 41565 28227 41568
rect 28169 41559 28227 41565
rect 28442 41556 28448 41568
rect 28500 41596 28506 41608
rect 29089 41599 29147 41605
rect 29089 41596 29101 41599
rect 28500 41568 29101 41596
rect 28500 41556 28506 41568
rect 29089 41565 29101 41568
rect 29135 41565 29147 41599
rect 29089 41559 29147 41565
rect 29178 41556 29184 41608
rect 29236 41556 29242 41608
rect 29288 41568 31754 41596
rect 25924 41500 26280 41528
rect 25924 41488 25930 41500
rect 27706 41488 27712 41540
rect 27764 41528 27770 41540
rect 29288 41528 29316 41568
rect 27764 41500 29316 41528
rect 27764 41488 27770 41500
rect 30374 41488 30380 41540
rect 30432 41528 30438 41540
rect 31570 41528 31576 41540
rect 30432 41500 31576 41528
rect 30432 41488 30438 41500
rect 31570 41488 31576 41500
rect 31628 41488 31634 41540
rect 31726 41528 31754 41568
rect 31938 41556 31944 41608
rect 31996 41556 32002 41608
rect 33870 41556 33876 41608
rect 33928 41596 33934 41608
rect 34241 41599 34299 41605
rect 34241 41596 34253 41599
rect 33928 41568 34253 41596
rect 33928 41556 33934 41568
rect 34241 41565 34253 41568
rect 34287 41565 34299 41599
rect 34241 41559 34299 41565
rect 36538 41556 36544 41608
rect 36596 41556 36602 41608
rect 37016 41605 37044 41636
rect 38378 41624 38384 41636
rect 38436 41624 38442 41676
rect 39592 41673 39620 41704
rect 43257 41701 43269 41735
rect 43303 41732 43315 41735
rect 43346 41732 43352 41744
rect 43303 41704 43352 41732
rect 43303 41701 43315 41704
rect 43257 41695 43315 41701
rect 43346 41692 43352 41704
rect 43404 41692 43410 41744
rect 44560 41732 44588 41772
rect 44729 41769 44741 41803
rect 44775 41800 44787 41803
rect 46382 41800 46388 41812
rect 44775 41772 46388 41800
rect 44775 41769 44787 41772
rect 44729 41763 44787 41769
rect 46382 41760 46388 41772
rect 46440 41760 46446 41812
rect 47026 41760 47032 41812
rect 47084 41760 47090 41812
rect 47210 41760 47216 41812
rect 47268 41800 47274 41812
rect 48961 41803 49019 41809
rect 48961 41800 48973 41803
rect 47268 41772 48973 41800
rect 47268 41760 47274 41772
rect 48961 41769 48973 41772
rect 49007 41769 49019 41803
rect 48961 41763 49019 41769
rect 49050 41760 49056 41812
rect 49108 41760 49114 41812
rect 49421 41803 49479 41809
rect 49421 41769 49433 41803
rect 49467 41800 49479 41803
rect 49510 41800 49516 41812
rect 49467 41772 49516 41800
rect 49467 41769 49479 41772
rect 49421 41763 49479 41769
rect 49510 41760 49516 41772
rect 49568 41760 49574 41812
rect 50246 41760 50252 41812
rect 50304 41760 50310 41812
rect 50617 41803 50675 41809
rect 50617 41769 50629 41803
rect 50663 41800 50675 41803
rect 51534 41800 51540 41812
rect 50663 41772 51540 41800
rect 50663 41769 50675 41772
rect 50617 41763 50675 41769
rect 51534 41760 51540 41772
rect 51592 41760 51598 41812
rect 51810 41760 51816 41812
rect 51868 41800 51874 41812
rect 53466 41800 53472 41812
rect 51868 41772 53472 41800
rect 51868 41760 51874 41772
rect 53466 41760 53472 41772
rect 53524 41800 53530 41812
rect 58342 41800 58348 41812
rect 53524 41772 58348 41800
rect 53524 41760 53530 41772
rect 45462 41732 45468 41744
rect 44560 41704 45468 41732
rect 45462 41692 45468 41704
rect 45520 41692 45526 41744
rect 46014 41692 46020 41744
rect 46072 41692 46078 41744
rect 46842 41692 46848 41744
rect 46900 41732 46906 41744
rect 47486 41732 47492 41744
rect 46900 41704 47492 41732
rect 46900 41692 46906 41704
rect 47486 41692 47492 41704
rect 47544 41692 47550 41744
rect 47854 41692 47860 41744
rect 47912 41732 47918 41744
rect 48317 41735 48375 41741
rect 48317 41732 48329 41735
rect 47912 41704 48329 41732
rect 47912 41692 47918 41704
rect 48317 41701 48329 41704
rect 48363 41701 48375 41735
rect 48317 41695 48375 41701
rect 50709 41735 50767 41741
rect 50709 41701 50721 41735
rect 50755 41732 50767 41735
rect 51442 41732 51448 41744
rect 50755 41704 51448 41732
rect 50755 41701 50767 41704
rect 50709 41695 50767 41701
rect 51442 41692 51448 41704
rect 51500 41692 51506 41744
rect 52454 41692 52460 41744
rect 52512 41692 52518 41744
rect 54128 41741 54156 41772
rect 58342 41760 58348 41772
rect 58400 41760 58406 41812
rect 54113 41735 54171 41741
rect 54113 41701 54125 41735
rect 54159 41701 54171 41735
rect 54113 41695 54171 41701
rect 39577 41667 39635 41673
rect 39577 41633 39589 41667
rect 39623 41633 39635 41667
rect 41322 41664 41328 41676
rect 40986 41636 41328 41664
rect 39577 41627 39635 41633
rect 41322 41624 41328 41636
rect 41380 41624 41386 41676
rect 44390 41636 44496 41664
rect 44468 41608 44496 41636
rect 45094 41624 45100 41676
rect 45152 41624 45158 41676
rect 47397 41667 47455 41673
rect 47397 41664 47409 41667
rect 46860 41636 47409 41664
rect 37001 41599 37059 41605
rect 37001 41565 37013 41599
rect 37047 41565 37059 41599
rect 37001 41559 37059 41565
rect 37093 41599 37151 41605
rect 37093 41565 37105 41599
rect 37139 41596 37151 41599
rect 37826 41596 37832 41608
rect 37139 41568 37832 41596
rect 37139 41565 37151 41568
rect 37093 41559 37151 41565
rect 37826 41556 37832 41568
rect 37884 41556 37890 41608
rect 39850 41556 39856 41608
rect 39908 41556 39914 41608
rect 40402 41556 40408 41608
rect 40460 41596 40466 41608
rect 42521 41599 42579 41605
rect 42521 41596 42533 41599
rect 40460 41568 42533 41596
rect 40460 41556 40466 41568
rect 42521 41565 42533 41568
rect 42567 41565 42579 41599
rect 42521 41559 42579 41565
rect 42702 41556 42708 41608
rect 42760 41556 42766 41608
rect 42794 41556 42800 41608
rect 42852 41596 42858 41608
rect 42981 41599 43039 41605
rect 42981 41596 42993 41599
rect 42852 41568 42993 41596
rect 42852 41556 42858 41568
rect 42981 41565 42993 41568
rect 43027 41596 43039 41599
rect 43346 41596 43352 41608
rect 43027 41568 43352 41596
rect 43027 41565 43039 41568
rect 42981 41559 43039 41565
rect 43346 41556 43352 41568
rect 43404 41556 43410 41608
rect 44450 41556 44456 41608
rect 44508 41556 44514 41608
rect 46860 41605 46888 41636
rect 47397 41633 47409 41636
rect 47443 41664 47455 41667
rect 47946 41664 47952 41676
rect 47443 41636 47952 41664
rect 47443 41633 47455 41636
rect 47397 41627 47455 41633
rect 47946 41624 47952 41636
rect 48004 41624 48010 41676
rect 48225 41667 48283 41673
rect 48225 41633 48237 41667
rect 48271 41664 48283 41667
rect 48590 41664 48596 41676
rect 48271 41636 48596 41664
rect 48271 41633 48283 41636
rect 48225 41627 48283 41633
rect 48590 41624 48596 41636
rect 48648 41624 48654 41676
rect 51077 41667 51135 41673
rect 51077 41633 51089 41667
rect 51123 41664 51135 41667
rect 51350 41664 51356 41676
rect 51123 41636 51356 41664
rect 51123 41633 51135 41636
rect 51077 41627 51135 41633
rect 51350 41624 51356 41636
rect 51408 41624 51414 41676
rect 54481 41667 54539 41673
rect 54481 41664 54493 41667
rect 53590 41636 54493 41664
rect 54481 41633 54493 41636
rect 54527 41664 54539 41667
rect 55122 41664 55128 41676
rect 54527 41636 55128 41664
rect 54527 41633 54539 41636
rect 54481 41627 54539 41633
rect 55122 41624 55128 41636
rect 55180 41624 55186 41676
rect 57698 41624 57704 41676
rect 57756 41624 57762 41676
rect 45373 41599 45431 41605
rect 45373 41565 45385 41599
rect 45419 41596 45431 41599
rect 46845 41599 46903 41605
rect 45419 41568 46520 41596
rect 45419 41565 45431 41568
rect 45373 41559 45431 41565
rect 31846 41528 31852 41540
rect 31726 41500 31852 41528
rect 31846 41488 31852 41500
rect 31904 41488 31910 41540
rect 33502 41488 33508 41540
rect 33560 41528 33566 41540
rect 34422 41528 34428 41540
rect 33560 41500 34428 41528
rect 33560 41488 33566 41500
rect 34422 41488 34428 41500
rect 34480 41528 34486 41540
rect 35253 41531 35311 41537
rect 35253 41528 35265 41531
rect 34480 41500 35265 41528
rect 34480 41488 34486 41500
rect 35253 41497 35265 41500
rect 35299 41497 35311 41531
rect 46492 41528 46520 41568
rect 46845 41565 46857 41599
rect 46891 41565 46903 41599
rect 46845 41559 46903 41565
rect 47578 41556 47584 41608
rect 47636 41556 47642 41608
rect 48409 41599 48467 41605
rect 48409 41565 48421 41599
rect 48455 41565 48467 41599
rect 48777 41599 48835 41605
rect 48777 41596 48789 41599
rect 48409 41559 48467 41565
rect 48516 41568 48789 41596
rect 47857 41531 47915 41537
rect 47857 41528 47869 41531
rect 46492 41500 47869 41528
rect 35253 41491 35311 41497
rect 47857 41497 47869 41500
rect 47903 41497 47915 41531
rect 47857 41491 47915 41497
rect 48222 41488 48228 41540
rect 48280 41528 48286 41540
rect 48424 41528 48452 41559
rect 48280 41500 48452 41528
rect 48280 41488 48286 41500
rect 21726 41460 21732 41472
rect 20732 41432 21732 41460
rect 20349 41423 20407 41429
rect 21726 41420 21732 41432
rect 21784 41420 21790 41472
rect 23106 41420 23112 41472
rect 23164 41460 23170 41472
rect 30466 41460 30472 41472
rect 23164 41432 30472 41460
rect 23164 41420 23170 41432
rect 30466 41420 30472 41432
rect 30524 41420 30530 41472
rect 30650 41420 30656 41472
rect 30708 41460 30714 41472
rect 32030 41460 32036 41472
rect 30708 41432 32036 41460
rect 30708 41420 30714 41432
rect 32030 41420 32036 41432
rect 32088 41420 32094 41472
rect 32398 41420 32404 41472
rect 32456 41460 32462 41472
rect 34514 41460 34520 41472
rect 32456 41432 34520 41460
rect 32456 41420 32462 41432
rect 34514 41420 34520 41432
rect 34572 41420 34578 41472
rect 34882 41420 34888 41472
rect 34940 41420 34946 41472
rect 35894 41420 35900 41472
rect 35952 41420 35958 41472
rect 37550 41420 37556 41472
rect 37608 41420 37614 41472
rect 41690 41420 41696 41472
rect 41748 41460 41754 41472
rect 42061 41463 42119 41469
rect 42061 41460 42073 41463
rect 41748 41432 42073 41460
rect 41748 41420 41754 41432
rect 42061 41429 42073 41432
rect 42107 41429 42119 41463
rect 42061 41423 42119 41429
rect 47762 41420 47768 41472
rect 47820 41460 47826 41472
rect 48516 41460 48544 41568
rect 48777 41565 48789 41568
rect 48823 41565 48835 41599
rect 48777 41559 48835 41565
rect 50798 41556 50804 41608
rect 50856 41556 50862 41608
rect 52181 41599 52239 41605
rect 52181 41596 52193 41599
rect 51046 41568 52193 41596
rect 49970 41488 49976 41540
rect 50028 41528 50034 41540
rect 50890 41528 50896 41540
rect 50028 41500 50896 41528
rect 50028 41488 50034 41500
rect 50890 41488 50896 41500
rect 50948 41528 50954 41540
rect 51046 41528 51074 41568
rect 52181 41565 52193 41568
rect 52227 41565 52239 41599
rect 52181 41559 52239 41565
rect 56134 41556 56140 41608
rect 56192 41556 56198 41608
rect 56413 41599 56471 41605
rect 56413 41565 56425 41599
rect 56459 41596 56471 41599
rect 56502 41596 56508 41608
rect 56459 41568 56508 41596
rect 56459 41565 56471 41568
rect 56413 41559 56471 41565
rect 56502 41556 56508 41568
rect 56560 41556 56566 41608
rect 57057 41599 57115 41605
rect 57057 41565 57069 41599
rect 57103 41565 57115 41599
rect 57057 41559 57115 41565
rect 50948 41500 51074 41528
rect 53929 41531 53987 41537
rect 50948 41488 50954 41500
rect 53929 41497 53941 41531
rect 53975 41528 53987 41531
rect 54110 41528 54116 41540
rect 53975 41500 54116 41528
rect 53975 41497 53987 41500
rect 53929 41491 53987 41497
rect 54110 41488 54116 41500
rect 54168 41528 54174 41540
rect 54938 41528 54944 41540
rect 54168 41500 54944 41528
rect 54168 41488 54174 41500
rect 54938 41488 54944 41500
rect 54996 41488 55002 41540
rect 57072 41528 57100 41559
rect 56336 41500 57100 41528
rect 47820 41432 48544 41460
rect 54665 41463 54723 41469
rect 47820 41420 47826 41432
rect 54665 41429 54677 41463
rect 54711 41460 54723 41463
rect 55674 41460 55680 41472
rect 54711 41432 55680 41460
rect 54711 41429 54723 41432
rect 54665 41423 54723 41429
rect 55674 41420 55680 41432
rect 55732 41460 55738 41472
rect 56336 41460 56364 41500
rect 55732 41432 56364 41460
rect 55732 41420 55738 41432
rect 56410 41420 56416 41472
rect 56468 41460 56474 41472
rect 56505 41463 56563 41469
rect 56505 41460 56517 41463
rect 56468 41432 56517 41460
rect 56468 41420 56474 41432
rect 56505 41429 56517 41432
rect 56551 41429 56563 41463
rect 56505 41423 56563 41429
rect 57609 41463 57667 41469
rect 57609 41429 57621 41463
rect 57655 41460 57667 41463
rect 57790 41460 57796 41472
rect 57655 41432 57796 41460
rect 57655 41429 57667 41432
rect 57609 41423 57667 41429
rect 57790 41420 57796 41432
rect 57848 41420 57854 41472
rect 552 41370 66424 41392
rect 552 41318 1998 41370
rect 2050 41318 2062 41370
rect 2114 41318 2126 41370
rect 2178 41318 2190 41370
rect 2242 41318 2254 41370
rect 2306 41318 50998 41370
rect 51050 41318 51062 41370
rect 51114 41318 51126 41370
rect 51178 41318 51190 41370
rect 51242 41318 51254 41370
rect 51306 41318 66424 41370
rect 552 41296 66424 41318
rect 13722 41216 13728 41268
rect 13780 41256 13786 41268
rect 15654 41256 15660 41268
rect 13780 41228 15660 41256
rect 13780 41216 13786 41228
rect 15654 41216 15660 41228
rect 15712 41216 15718 41268
rect 16758 41216 16764 41268
rect 16816 41216 16822 41268
rect 19889 41259 19947 41265
rect 19889 41225 19901 41259
rect 19935 41256 19947 41259
rect 20990 41256 20996 41268
rect 19935 41228 20996 41256
rect 19935 41225 19947 41228
rect 19889 41219 19947 41225
rect 20990 41216 20996 41228
rect 21048 41216 21054 41268
rect 21542 41216 21548 41268
rect 21600 41256 21606 41268
rect 21821 41259 21879 41265
rect 21821 41256 21833 41259
rect 21600 41228 21833 41256
rect 21600 41216 21606 41228
rect 21821 41225 21833 41228
rect 21867 41225 21879 41259
rect 21821 41219 21879 41225
rect 23750 41216 23756 41268
rect 23808 41256 23814 41268
rect 24121 41259 24179 41265
rect 24121 41256 24133 41259
rect 23808 41228 24133 41256
rect 23808 41216 23814 41228
rect 24121 41225 24133 41228
rect 24167 41225 24179 41259
rect 25590 41256 25596 41268
rect 24121 41219 24179 41225
rect 24412 41228 25596 41256
rect 13078 41148 13084 41200
rect 13136 41188 13142 41200
rect 14642 41188 14648 41200
rect 13136 41160 14648 41188
rect 13136 41148 13142 41160
rect 8754 41080 8760 41132
rect 8812 41120 8818 41132
rect 9401 41123 9459 41129
rect 9401 41120 9413 41123
rect 8812 41092 9413 41120
rect 8812 41080 8818 41092
rect 9401 41089 9413 41092
rect 9447 41089 9459 41123
rect 9401 41083 9459 41089
rect 9677 41123 9735 41129
rect 9677 41089 9689 41123
rect 9723 41120 9735 41123
rect 10042 41120 10048 41132
rect 9723 41092 10048 41120
rect 9723 41089 9735 41092
rect 9677 41083 9735 41089
rect 10042 41080 10048 41092
rect 10100 41080 10106 41132
rect 11422 41080 11428 41132
rect 11480 41080 11486 41132
rect 11609 41123 11667 41129
rect 11609 41089 11621 41123
rect 11655 41120 11667 41123
rect 12434 41120 12440 41132
rect 11655 41092 12440 41120
rect 11655 41089 11667 41092
rect 11609 41083 11667 41089
rect 12434 41080 12440 41092
rect 12492 41080 12498 41132
rect 13740 41129 13768 41160
rect 14642 41148 14648 41160
rect 14700 41148 14706 41200
rect 19150 41188 19156 41200
rect 16316 41160 19156 41188
rect 13357 41123 13415 41129
rect 13357 41089 13369 41123
rect 13403 41089 13415 41123
rect 13357 41083 13415 41089
rect 13725 41123 13783 41129
rect 13725 41089 13737 41123
rect 13771 41089 13783 41123
rect 16316 41120 16344 41160
rect 19150 41148 19156 41160
rect 19208 41148 19214 41200
rect 21726 41148 21732 41200
rect 21784 41188 21790 41200
rect 22554 41188 22560 41200
rect 21784 41160 22560 41188
rect 21784 41148 21790 41160
rect 22554 41148 22560 41160
rect 22612 41148 22618 41200
rect 13725 41083 13783 41089
rect 14108 41092 16344 41120
rect 9309 41055 9367 41061
rect 9309 41021 9321 41055
rect 9355 41021 9367 41055
rect 13372 41052 13400 41083
rect 13814 41052 13820 41064
rect 13372 41024 13820 41052
rect 9309 41015 9367 41021
rect 9324 40984 9352 41015
rect 13814 41012 13820 41024
rect 13872 41052 13878 41064
rect 13909 41055 13967 41061
rect 13909 41052 13921 41055
rect 13872 41024 13921 41052
rect 13872 41012 13878 41024
rect 13909 41021 13921 41024
rect 13955 41021 13967 41055
rect 13909 41015 13967 41021
rect 9674 40984 9680 40996
rect 9324 40956 9680 40984
rect 9674 40944 9680 40956
rect 9732 40944 9738 40996
rect 9766 40944 9772 40996
rect 9824 40984 9830 40996
rect 10134 40984 10140 40996
rect 9824 40956 10140 40984
rect 9824 40944 9830 40956
rect 10134 40944 10140 40956
rect 10192 40944 10198 40996
rect 11882 40944 11888 40996
rect 11940 40944 11946 40996
rect 12894 40944 12900 40996
rect 12952 40944 12958 40996
rect 14108 40984 14136 41092
rect 17494 41080 17500 41132
rect 17552 41120 17558 41132
rect 17862 41120 17868 41132
rect 17552 41092 17868 41120
rect 17552 41080 17558 41092
rect 17862 41080 17868 41092
rect 17920 41080 17926 41132
rect 17954 41080 17960 41132
rect 18012 41120 18018 41132
rect 18417 41123 18475 41129
rect 18417 41120 18429 41123
rect 18012 41092 18429 41120
rect 18012 41080 18018 41092
rect 18417 41089 18429 41092
rect 18463 41089 18475 41123
rect 18417 41083 18475 41089
rect 19978 41080 19984 41132
rect 20036 41080 20042 41132
rect 20254 41080 20260 41132
rect 20312 41080 20318 41132
rect 21450 41080 21456 41132
rect 21508 41120 21514 41132
rect 22373 41123 22431 41129
rect 22373 41120 22385 41123
rect 21508 41092 22385 41120
rect 21508 41080 21514 41092
rect 22373 41089 22385 41092
rect 22419 41089 22431 41123
rect 22373 41083 22431 41089
rect 23109 41123 23167 41129
rect 23109 41089 23121 41123
rect 23155 41120 23167 41123
rect 24412 41120 24440 41228
rect 25590 41216 25596 41228
rect 25648 41216 25654 41268
rect 25685 41259 25743 41265
rect 25685 41225 25697 41259
rect 25731 41256 25743 41259
rect 26234 41256 26240 41268
rect 25731 41228 26240 41256
rect 25731 41225 25743 41228
rect 25685 41219 25743 41225
rect 26234 41216 26240 41228
rect 26292 41256 26298 41268
rect 26970 41256 26976 41268
rect 26292 41228 26976 41256
rect 26292 41216 26298 41228
rect 26970 41216 26976 41228
rect 27028 41216 27034 41268
rect 27154 41216 27160 41268
rect 27212 41256 27218 41268
rect 27212 41228 33824 41256
rect 27212 41216 27218 41228
rect 25222 41148 25228 41200
rect 25280 41188 25286 41200
rect 25866 41188 25872 41200
rect 25280 41160 25872 41188
rect 25280 41148 25286 41160
rect 25866 41148 25872 41160
rect 25924 41148 25930 41200
rect 33796 41188 33824 41228
rect 33870 41216 33876 41268
rect 33928 41216 33934 41268
rect 35802 41256 35808 41268
rect 33980 41228 35808 41256
rect 33980 41188 34008 41228
rect 35802 41216 35808 41228
rect 35860 41216 35866 41268
rect 37090 41216 37096 41268
rect 37148 41256 37154 41268
rect 37645 41259 37703 41265
rect 37645 41256 37657 41259
rect 37148 41228 37657 41256
rect 37148 41216 37154 41228
rect 37645 41225 37657 41228
rect 37691 41225 37703 41259
rect 37645 41219 37703 41225
rect 37826 41216 37832 41268
rect 37884 41216 37890 41268
rect 39114 41216 39120 41268
rect 39172 41256 39178 41268
rect 39301 41259 39359 41265
rect 39301 41256 39313 41259
rect 39172 41228 39313 41256
rect 39172 41216 39178 41228
rect 39301 41225 39313 41228
rect 39347 41225 39359 41259
rect 39301 41219 39359 41225
rect 39482 41216 39488 41268
rect 39540 41256 39546 41268
rect 39540 41228 42748 41256
rect 39540 41216 39546 41228
rect 25976 41160 32076 41188
rect 33796 41160 34008 41188
rect 34149 41191 34207 41197
rect 24670 41120 24676 41132
rect 23155 41092 24440 41120
rect 24504 41092 24676 41120
rect 23155 41089 23167 41092
rect 23109 41083 23167 41089
rect 15013 41055 15071 41061
rect 15013 41021 15025 41055
rect 15059 41021 15071 41055
rect 15013 41015 15071 41021
rect 17221 41055 17279 41061
rect 17221 41021 17233 41055
rect 17267 41052 17279 41055
rect 18046 41052 18052 41064
rect 17267 41024 18052 41052
rect 17267 41021 17279 41024
rect 17221 41015 17279 41021
rect 13740 40956 14136 40984
rect 15028 40984 15056 41015
rect 18046 41012 18052 41024
rect 18104 41012 18110 41064
rect 19058 41012 19064 41064
rect 19116 41052 19122 41064
rect 19245 41055 19303 41061
rect 19245 41052 19257 41055
rect 19116 41024 19257 41052
rect 19116 41012 19122 41024
rect 19245 41021 19257 41024
rect 19291 41021 19303 41055
rect 19245 41015 19303 41021
rect 23014 41012 23020 41064
rect 23072 41052 23078 41064
rect 24504 41052 24532 41092
rect 24670 41080 24676 41092
rect 24728 41080 24734 41132
rect 25130 41080 25136 41132
rect 25188 41120 25194 41132
rect 25976 41120 26004 41160
rect 25188 41092 26004 41120
rect 25188 41080 25194 41092
rect 26878 41080 26884 41132
rect 26936 41120 26942 41132
rect 30469 41123 30527 41129
rect 26936 41092 27476 41120
rect 26936 41080 26942 41092
rect 27448 41064 27476 41092
rect 30469 41089 30481 41123
rect 30515 41120 30527 41123
rect 31110 41120 31116 41132
rect 30515 41092 31116 41120
rect 30515 41089 30527 41092
rect 30469 41083 30527 41089
rect 31110 41080 31116 41092
rect 31168 41080 31174 41132
rect 31570 41080 31576 41132
rect 31628 41120 31634 41132
rect 31849 41123 31907 41129
rect 31849 41120 31861 41123
rect 31628 41092 31861 41120
rect 31628 41080 31634 41092
rect 31849 41089 31861 41092
rect 31895 41089 31907 41123
rect 31849 41083 31907 41089
rect 23072 41024 24532 41052
rect 24581 41055 24639 41061
rect 23072 41012 23078 41024
rect 24581 41021 24593 41055
rect 24627 41052 24639 41055
rect 24762 41052 24768 41064
rect 24627 41024 24768 41052
rect 24627 41021 24639 41024
rect 24581 41015 24639 41021
rect 24762 41012 24768 41024
rect 24820 41012 24826 41064
rect 26973 41055 27031 41061
rect 26973 41052 26985 41055
rect 25240 41024 26985 41052
rect 15194 40984 15200 40996
rect 15028 40956 15200 40984
rect 8665 40919 8723 40925
rect 8665 40885 8677 40919
rect 8711 40916 8723 40919
rect 8938 40916 8944 40928
rect 8711 40888 8944 40916
rect 8711 40885 8723 40888
rect 8665 40879 8723 40885
rect 8938 40876 8944 40888
rect 8996 40876 9002 40928
rect 11422 40876 11428 40928
rect 11480 40916 11486 40928
rect 12802 40916 12808 40928
rect 11480 40888 12808 40916
rect 11480 40876 11486 40888
rect 12802 40876 12808 40888
rect 12860 40916 12866 40928
rect 13740 40916 13768 40956
rect 15194 40944 15200 40956
rect 15252 40944 15258 40996
rect 15286 40944 15292 40996
rect 15344 40944 15350 40996
rect 16298 40944 16304 40996
rect 16356 40944 16362 40996
rect 18782 40944 18788 40996
rect 18840 40984 18846 40996
rect 18840 40956 20024 40984
rect 18840 40944 18846 40956
rect 12860 40888 13768 40916
rect 12860 40876 12866 40888
rect 13814 40876 13820 40928
rect 13872 40876 13878 40928
rect 14090 40876 14096 40928
rect 14148 40916 14154 40928
rect 14277 40919 14335 40925
rect 14277 40916 14289 40919
rect 14148 40888 14289 40916
rect 14148 40876 14154 40888
rect 14277 40885 14289 40888
rect 14323 40885 14335 40919
rect 14277 40879 14335 40885
rect 14458 40876 14464 40928
rect 14516 40916 14522 40928
rect 16853 40919 16911 40925
rect 16853 40916 16865 40919
rect 14516 40888 16865 40916
rect 14516 40876 14522 40888
rect 16853 40885 16865 40888
rect 16899 40885 16911 40919
rect 16853 40879 16911 40885
rect 16942 40876 16948 40928
rect 17000 40916 17006 40928
rect 17313 40919 17371 40925
rect 17313 40916 17325 40919
rect 17000 40888 17325 40916
rect 17000 40876 17006 40888
rect 17313 40885 17325 40888
rect 17359 40885 17371 40919
rect 17313 40879 17371 40885
rect 17402 40876 17408 40928
rect 17460 40916 17466 40928
rect 17865 40919 17923 40925
rect 17865 40916 17877 40919
rect 17460 40888 17877 40916
rect 17460 40876 17466 40888
rect 17865 40885 17877 40888
rect 17911 40885 17923 40919
rect 19996 40916 20024 40956
rect 20346 40944 20352 40996
rect 20404 40984 20410 40996
rect 25240 40984 25268 41024
rect 26973 41021 26985 41024
rect 27019 41021 27031 41055
rect 26973 41015 27031 41021
rect 20404 40956 20746 40984
rect 21560 40956 25268 40984
rect 26988 40984 27016 41015
rect 27062 41012 27068 41064
rect 27120 41012 27126 41064
rect 27430 41012 27436 41064
rect 27488 41052 27494 41064
rect 28813 41055 28871 41061
rect 28813 41052 28825 41055
rect 27488 41024 28825 41052
rect 27488 41012 27494 41024
rect 28813 41021 28825 41024
rect 28859 41052 28871 41055
rect 30098 41052 30104 41064
rect 28859 41024 30104 41052
rect 28859 41021 28871 41024
rect 28813 41015 28871 41021
rect 30098 41012 30104 41024
rect 30156 41012 30162 41064
rect 30650 41012 30656 41064
rect 30708 41012 30714 41064
rect 31205 41055 31263 41061
rect 31205 41021 31217 41055
rect 31251 41052 31263 41055
rect 31665 41055 31723 41061
rect 31665 41052 31677 41055
rect 31251 41024 31677 41052
rect 31251 41021 31263 41024
rect 31205 41015 31263 41021
rect 31665 41021 31677 41024
rect 31711 41021 31723 41055
rect 32048 41052 32076 41160
rect 34149 41157 34161 41191
rect 34195 41157 34207 41191
rect 34149 41151 34207 41157
rect 32122 41080 32128 41132
rect 32180 41080 32186 41132
rect 32401 41123 32459 41129
rect 32401 41089 32413 41123
rect 32447 41120 32459 41123
rect 34164 41120 34192 41151
rect 32447 41092 34192 41120
rect 32447 41089 32459 41092
rect 32401 41083 32459 41089
rect 34238 41080 34244 41132
rect 34296 41120 34302 41132
rect 34701 41123 34759 41129
rect 34701 41120 34713 41123
rect 34296 41092 34713 41120
rect 34296 41080 34302 41092
rect 34701 41089 34713 41092
rect 34747 41089 34759 41123
rect 34701 41083 34759 41089
rect 35250 41080 35256 41132
rect 35308 41120 35314 41132
rect 35529 41123 35587 41129
rect 35529 41120 35541 41123
rect 35308 41092 35541 41120
rect 35308 41080 35314 41092
rect 35529 41089 35541 41092
rect 35575 41120 35587 41123
rect 35710 41120 35716 41132
rect 35575 41092 35716 41120
rect 35575 41089 35587 41092
rect 35529 41083 35587 41089
rect 35710 41080 35716 41092
rect 35768 41080 35774 41132
rect 35894 41080 35900 41132
rect 35952 41080 35958 41132
rect 34517 41055 34575 41061
rect 32048 41024 32168 41052
rect 31665 41015 31723 41021
rect 31846 40984 31852 40996
rect 26988 40956 31852 40984
rect 20404 40944 20410 40956
rect 21560 40916 21588 40956
rect 31846 40944 31852 40956
rect 31904 40944 31910 40996
rect 32140 40984 32168 41024
rect 34517 41021 34529 41055
rect 34563 41052 34575 41055
rect 34882 41052 34888 41064
rect 34563 41024 34888 41052
rect 34563 41021 34575 41024
rect 34517 41015 34575 41021
rect 34882 41012 34888 41024
rect 34940 41012 34946 41064
rect 35345 41055 35403 41061
rect 35345 41021 35357 41055
rect 35391 41052 35403 41055
rect 35912 41052 35940 41080
rect 37108 41052 37136 41216
rect 42720 41200 42748 41228
rect 47854 41216 47860 41268
rect 47912 41216 47918 41268
rect 48590 41216 48596 41268
rect 48648 41216 48654 41268
rect 52270 41216 52276 41268
rect 52328 41256 52334 41268
rect 53009 41259 53067 41265
rect 52328 41228 52684 41256
rect 52328 41216 52334 41228
rect 38930 41188 38936 41200
rect 38304 41160 38936 41188
rect 38304 41129 38332 41160
rect 38930 41148 38936 41160
rect 38988 41148 38994 41200
rect 40126 41188 40132 41200
rect 39684 41160 40132 41188
rect 38289 41123 38347 41129
rect 38289 41089 38301 41123
rect 38335 41089 38347 41123
rect 38289 41083 38347 41089
rect 38473 41123 38531 41129
rect 38473 41089 38485 41123
rect 38519 41120 38531 41123
rect 39684 41120 39712 41160
rect 38519 41092 39712 41120
rect 38519 41089 38531 41092
rect 38473 41083 38531 41089
rect 39758 41080 39764 41132
rect 39816 41080 39822 41132
rect 39868 41129 39896 41160
rect 40126 41148 40132 41160
rect 40184 41188 40190 41200
rect 40678 41188 40684 41200
rect 40184 41160 40684 41188
rect 40184 41148 40190 41160
rect 40678 41148 40684 41160
rect 40736 41148 40742 41200
rect 42702 41148 42708 41200
rect 42760 41188 42766 41200
rect 42760 41160 43208 41188
rect 42760 41148 42766 41160
rect 39853 41123 39911 41129
rect 39853 41089 39865 41123
rect 39899 41089 39911 41123
rect 43070 41120 43076 41132
rect 39853 41083 39911 41089
rect 40420 41092 43076 41120
rect 35391 41024 35940 41052
rect 37016 41024 37136 41052
rect 35391 41021 35403 41024
rect 35345 41015 35403 41021
rect 34146 40984 34152 40996
rect 32140 40956 32352 40984
rect 33626 40956 34152 40984
rect 19996 40888 21588 40916
rect 17865 40879 17923 40885
rect 22186 40876 22192 40928
rect 22244 40876 22250 40928
rect 22278 40876 22284 40928
rect 22336 40876 22342 40928
rect 23661 40919 23719 40925
rect 23661 40885 23673 40919
rect 23707 40916 23719 40919
rect 24394 40916 24400 40928
rect 23707 40888 24400 40916
rect 23707 40885 23719 40888
rect 23661 40879 23719 40885
rect 24394 40876 24400 40888
rect 24452 40876 24458 40928
rect 24489 40919 24547 40925
rect 24489 40885 24501 40919
rect 24535 40916 24547 40919
rect 24670 40916 24676 40928
rect 24535 40888 24676 40916
rect 24535 40885 24547 40888
rect 24489 40879 24547 40885
rect 24670 40876 24676 40888
rect 24728 40876 24734 40928
rect 24854 40876 24860 40928
rect 24912 40916 24918 40928
rect 27522 40916 27528 40928
rect 24912 40888 27528 40916
rect 24912 40876 24918 40888
rect 27522 40876 27528 40888
rect 27580 40876 27586 40928
rect 29086 40876 29092 40928
rect 29144 40916 29150 40928
rect 29825 40919 29883 40925
rect 29825 40916 29837 40919
rect 29144 40888 29837 40916
rect 29144 40876 29150 40888
rect 29825 40885 29837 40888
rect 29871 40885 29883 40919
rect 29825 40879 29883 40885
rect 29914 40876 29920 40928
rect 29972 40916 29978 40928
rect 31297 40919 31355 40925
rect 31297 40916 31309 40919
rect 29972 40888 31309 40916
rect 29972 40876 29978 40888
rect 31297 40885 31309 40888
rect 31343 40885 31355 40919
rect 31297 40879 31355 40885
rect 31757 40919 31815 40925
rect 31757 40885 31769 40919
rect 31803 40916 31815 40919
rect 32214 40916 32220 40928
rect 31803 40888 32220 40916
rect 31803 40885 31815 40888
rect 31757 40879 31815 40885
rect 32214 40876 32220 40888
rect 32272 40876 32278 40928
rect 32324 40916 32352 40956
rect 34146 40944 34152 40956
rect 34204 40944 34210 40996
rect 35894 40944 35900 40996
rect 35952 40984 35958 40996
rect 36262 40984 36268 40996
rect 35952 40956 36268 40984
rect 35952 40944 35958 40956
rect 36262 40944 36268 40956
rect 36320 40944 36326 40996
rect 33410 40916 33416 40928
rect 32324 40888 33416 40916
rect 33410 40876 33416 40888
rect 33468 40876 33474 40928
rect 34606 40876 34612 40928
rect 34664 40876 34670 40928
rect 34977 40919 35035 40925
rect 34977 40885 34989 40919
rect 35023 40916 35035 40919
rect 35066 40916 35072 40928
rect 35023 40888 35072 40916
rect 35023 40885 35035 40888
rect 34977 40879 35035 40885
rect 35066 40876 35072 40888
rect 35124 40876 35130 40928
rect 35434 40876 35440 40928
rect 35492 40876 35498 40928
rect 37016 40916 37044 41024
rect 37182 41012 37188 41064
rect 37240 41052 37246 41064
rect 38657 41055 38715 41061
rect 38657 41052 38669 41055
rect 37240 41024 38669 41052
rect 37240 41012 37246 41024
rect 38657 41021 38669 41024
rect 38703 41021 38715 41055
rect 38657 41015 38715 41021
rect 37090 40944 37096 40996
rect 37148 40984 37154 40996
rect 37553 40987 37611 40993
rect 37553 40984 37565 40987
rect 37148 40956 37565 40984
rect 37148 40944 37154 40956
rect 37553 40953 37565 40956
rect 37599 40984 37611 40987
rect 40420 40984 40448 41092
rect 43070 41080 43076 41092
rect 43128 41080 43134 41132
rect 43180 41129 43208 41160
rect 46106 41148 46112 41200
rect 46164 41188 46170 41200
rect 52546 41188 52552 41200
rect 46164 41160 52552 41188
rect 46164 41148 46170 41160
rect 52546 41148 52552 41160
rect 52604 41148 52610 41200
rect 52656 41188 52684 41228
rect 53009 41225 53021 41259
rect 53055 41256 53067 41259
rect 53190 41256 53196 41268
rect 53055 41228 53196 41256
rect 53055 41225 53067 41228
rect 53009 41219 53067 41225
rect 53190 41216 53196 41228
rect 53248 41216 53254 41268
rect 57698 41256 57704 41268
rect 53300 41228 57704 41256
rect 53300 41188 53328 41228
rect 57698 41216 57704 41228
rect 57756 41216 57762 41268
rect 54018 41188 54024 41200
rect 52656 41160 53328 41188
rect 53484 41160 54024 41188
rect 43165 41123 43223 41129
rect 43165 41089 43177 41123
rect 43211 41120 43223 41123
rect 46937 41123 46995 41129
rect 43211 41092 43484 41120
rect 43211 41089 43223 41092
rect 43165 41083 43223 41089
rect 41966 41012 41972 41064
rect 42024 41052 42030 41064
rect 42794 41052 42800 41064
rect 42024 41024 42800 41052
rect 42024 41012 42030 41024
rect 42794 41012 42800 41024
rect 42852 41012 42858 41064
rect 43456 41052 43484 41092
rect 46937 41089 46949 41123
rect 46983 41089 46995 41123
rect 46937 41083 46995 41089
rect 47305 41123 47363 41129
rect 47305 41089 47317 41123
rect 47351 41120 47363 41123
rect 47854 41120 47860 41132
rect 47351 41092 47860 41120
rect 47351 41089 47363 41092
rect 47305 41083 47363 41089
rect 45002 41052 45008 41064
rect 43456 41024 45008 41052
rect 45002 41012 45008 41024
rect 45060 41052 45066 41064
rect 46952 41052 46980 41083
rect 47854 41080 47860 41092
rect 47912 41080 47918 41132
rect 47946 41080 47952 41132
rect 48004 41080 48010 41132
rect 48774 41080 48780 41132
rect 48832 41120 48838 41132
rect 49326 41120 49332 41132
rect 48832 41092 49332 41120
rect 48832 41080 48838 41092
rect 49326 41080 49332 41092
rect 49384 41120 49390 41132
rect 50249 41123 50307 41129
rect 50249 41120 50261 41123
rect 49384 41092 50261 41120
rect 49384 41080 49390 41092
rect 50249 41089 50261 41092
rect 50295 41089 50307 41123
rect 50249 41083 50307 41089
rect 50264 41052 50292 41083
rect 50614 41080 50620 41132
rect 50672 41120 50678 41132
rect 53484 41129 53512 41160
rect 54018 41148 54024 41160
rect 54076 41148 54082 41200
rect 54478 41188 54484 41200
rect 54128 41160 54484 41188
rect 53469 41123 53527 41129
rect 53469 41120 53481 41123
rect 50672 41092 53481 41120
rect 50672 41080 50678 41092
rect 53469 41089 53481 41092
rect 53515 41089 53527 41123
rect 53469 41083 53527 41089
rect 53650 41080 53656 41132
rect 53708 41080 53714 41132
rect 53929 41123 53987 41129
rect 53929 41089 53941 41123
rect 53975 41120 53987 41123
rect 54128 41120 54156 41160
rect 54478 41148 54484 41160
rect 54536 41148 54542 41200
rect 54846 41148 54852 41200
rect 54904 41188 54910 41200
rect 54904 41160 60734 41188
rect 54904 41148 54910 41160
rect 53975 41092 54156 41120
rect 53975 41089 53987 41092
rect 53929 41083 53987 41089
rect 54202 41080 54208 41132
rect 54260 41120 54266 41132
rect 55030 41120 55036 41132
rect 54260 41092 55036 41120
rect 54260 41080 54266 41092
rect 55030 41080 55036 41092
rect 55088 41120 55094 41132
rect 55861 41123 55919 41129
rect 55861 41120 55873 41123
rect 55088 41092 55873 41120
rect 55088 41080 55094 41092
rect 55861 41089 55873 41092
rect 55907 41089 55919 41123
rect 55861 41083 55919 41089
rect 55968 41092 56640 41120
rect 51074 41052 51080 41064
rect 45060 41024 50200 41052
rect 50264 41024 51080 41052
rect 45060 41012 45066 41024
rect 41414 40984 41420 40996
rect 37599 40956 40448 40984
rect 41262 40956 41420 40984
rect 37599 40953 37611 40956
rect 37553 40947 37611 40953
rect 41414 40944 41420 40956
rect 41472 40984 41478 40996
rect 41598 40984 41604 40996
rect 41472 40956 41604 40984
rect 41472 40944 41478 40956
rect 41598 40944 41604 40956
rect 41656 40944 41662 40996
rect 41690 40944 41696 40996
rect 41748 40944 41754 40996
rect 42242 40944 42248 40996
rect 42300 40984 42306 40996
rect 42981 40987 43039 40993
rect 42981 40984 42993 40987
rect 42300 40956 42993 40984
rect 42300 40944 42306 40956
rect 42981 40953 42993 40956
rect 43027 40953 43039 40987
rect 42981 40947 43039 40953
rect 43162 40944 43168 40996
rect 43220 40984 43226 40996
rect 43349 40987 43407 40993
rect 43349 40984 43361 40987
rect 43220 40956 43361 40984
rect 43220 40944 43226 40956
rect 43349 40953 43361 40956
rect 43395 40984 43407 40987
rect 44453 40987 44511 40993
rect 44453 40984 44465 40987
rect 43395 40956 44465 40984
rect 43395 40953 43407 40956
rect 43349 40947 43407 40953
rect 44453 40953 44465 40956
rect 44499 40984 44511 40987
rect 45094 40984 45100 40996
rect 44499 40956 45100 40984
rect 44499 40953 44511 40956
rect 44453 40947 44511 40953
rect 45094 40944 45100 40956
rect 45152 40984 45158 40996
rect 45462 40984 45468 40996
rect 45152 40956 45468 40984
rect 45152 40944 45158 40956
rect 45462 40944 45468 40956
rect 45520 40944 45526 40996
rect 46201 40987 46259 40993
rect 46201 40953 46213 40987
rect 46247 40953 46259 40987
rect 46201 40947 46259 40953
rect 38197 40919 38255 40925
rect 38197 40916 38209 40919
rect 37016 40888 38209 40916
rect 38197 40885 38209 40888
rect 38243 40885 38255 40919
rect 38197 40879 38255 40885
rect 39669 40919 39727 40925
rect 39669 40885 39681 40919
rect 39715 40916 39727 40919
rect 40034 40916 40040 40928
rect 39715 40888 40040 40916
rect 39715 40885 39727 40888
rect 39669 40879 39727 40885
rect 40034 40876 40040 40888
rect 40092 40876 40098 40928
rect 40221 40919 40279 40925
rect 40221 40885 40233 40919
rect 40267 40916 40279 40919
rect 40402 40916 40408 40928
rect 40267 40888 40408 40916
rect 40267 40885 40279 40888
rect 40221 40879 40279 40885
rect 40402 40876 40408 40888
rect 40460 40916 40466 40928
rect 40954 40916 40960 40928
rect 40460 40888 40960 40916
rect 40460 40876 40466 40888
rect 40954 40876 40960 40888
rect 41012 40876 41018 40928
rect 42521 40919 42579 40925
rect 42521 40885 42533 40919
rect 42567 40916 42579 40919
rect 42794 40916 42800 40928
rect 42567 40888 42800 40916
rect 42567 40885 42579 40888
rect 42521 40879 42579 40885
rect 42794 40876 42800 40888
rect 42852 40876 42858 40928
rect 42886 40876 42892 40928
rect 42944 40876 42950 40928
rect 43070 40876 43076 40928
rect 43128 40916 43134 40928
rect 46106 40916 46112 40928
rect 43128 40888 46112 40916
rect 43128 40876 43134 40888
rect 46106 40876 46112 40888
rect 46164 40916 46170 40928
rect 46216 40916 46244 40947
rect 46474 40944 46480 40996
rect 46532 40984 46538 40996
rect 46753 40987 46811 40993
rect 46753 40984 46765 40987
rect 46532 40956 46765 40984
rect 46532 40944 46538 40956
rect 46753 40953 46765 40956
rect 46799 40984 46811 40987
rect 47397 40987 47455 40993
rect 47397 40984 47409 40987
rect 46799 40956 47409 40984
rect 46799 40953 46811 40956
rect 46753 40947 46811 40953
rect 47397 40953 47409 40956
rect 47443 40953 47455 40987
rect 47397 40947 47455 40953
rect 47486 40944 47492 40996
rect 47544 40944 47550 40996
rect 48038 40944 48044 40996
rect 48096 40984 48102 40996
rect 49510 40984 49516 40996
rect 48096 40956 49516 40984
rect 48096 40944 48102 40956
rect 49510 40944 49516 40956
rect 49568 40944 49574 40996
rect 49602 40944 49608 40996
rect 49660 40984 49666 40996
rect 50065 40987 50123 40993
rect 50065 40984 50077 40987
rect 49660 40956 50077 40984
rect 49660 40944 49666 40956
rect 50065 40953 50077 40956
rect 50111 40953 50123 40987
rect 50172 40984 50200 41024
rect 51074 41012 51080 41024
rect 51132 41012 51138 41064
rect 51166 41012 51172 41064
rect 51224 41052 51230 41064
rect 55968 41052 55996 41092
rect 51224 41024 55996 41052
rect 51224 41012 51230 41024
rect 56410 41012 56416 41064
rect 56468 41052 56474 41064
rect 56505 41055 56563 41061
rect 56505 41052 56517 41055
rect 56468 41024 56517 41052
rect 56468 41012 56474 41024
rect 56505 41021 56517 41024
rect 56551 41021 56563 41055
rect 56612 41052 56640 41092
rect 56686 41080 56692 41132
rect 56744 41080 56750 41132
rect 57054 41080 57060 41132
rect 57112 41120 57118 41132
rect 57517 41123 57575 41129
rect 57517 41120 57529 41123
rect 57112 41092 57529 41120
rect 57112 41080 57118 41092
rect 57517 41089 57529 41092
rect 57563 41089 57575 41123
rect 57517 41083 57575 41089
rect 56612 41024 57284 41052
rect 56505 41015 56563 41021
rect 54205 40987 54263 40993
rect 50172 40956 54156 40984
rect 50065 40947 50123 40953
rect 46164 40888 46244 40916
rect 46164 40876 46170 40888
rect 46290 40876 46296 40928
rect 46348 40876 46354 40928
rect 46658 40876 46664 40928
rect 46716 40876 46722 40928
rect 49418 40876 49424 40928
rect 49476 40916 49482 40928
rect 49697 40919 49755 40925
rect 49697 40916 49709 40919
rect 49476 40888 49709 40916
rect 49476 40876 49482 40888
rect 49697 40885 49709 40888
rect 49743 40885 49755 40919
rect 49697 40879 49755 40885
rect 50154 40876 50160 40928
rect 50212 40876 50218 40928
rect 51350 40876 51356 40928
rect 51408 40916 51414 40928
rect 52362 40916 52368 40928
rect 51408 40888 52368 40916
rect 51408 40876 51414 40888
rect 52362 40876 52368 40888
rect 52420 40916 52426 40928
rect 52457 40919 52515 40925
rect 52457 40916 52469 40919
rect 52420 40888 52469 40916
rect 52420 40876 52426 40888
rect 52457 40885 52469 40888
rect 52503 40885 52515 40919
rect 52457 40879 52515 40885
rect 52822 40876 52828 40928
rect 52880 40916 52886 40928
rect 53377 40919 53435 40925
rect 53377 40916 53389 40919
rect 52880 40888 53389 40916
rect 52880 40876 52886 40888
rect 53377 40885 53389 40888
rect 53423 40885 53435 40919
rect 54128 40916 54156 40956
rect 54205 40953 54217 40987
rect 54251 40984 54263 40987
rect 54754 40984 54760 40996
rect 54251 40956 54760 40984
rect 54251 40953 54263 40956
rect 54205 40947 54263 40953
rect 54754 40944 54760 40956
rect 54812 40944 54818 40996
rect 54849 40987 54907 40993
rect 54849 40953 54861 40987
rect 54895 40984 54907 40987
rect 54895 40956 56364 40984
rect 54895 40953 54907 40956
rect 54849 40947 54907 40953
rect 54864 40916 54892 40947
rect 54128 40888 54892 40916
rect 54941 40919 54999 40925
rect 53377 40879 53435 40885
rect 54941 40885 54953 40919
rect 54987 40916 54999 40919
rect 55030 40916 55036 40928
rect 54987 40888 55036 40916
rect 54987 40885 54999 40888
rect 54941 40879 54999 40885
rect 55030 40876 55036 40888
rect 55088 40876 55094 40928
rect 55214 40876 55220 40928
rect 55272 40916 55278 40928
rect 55309 40919 55367 40925
rect 55309 40916 55321 40919
rect 55272 40888 55321 40916
rect 55272 40876 55278 40888
rect 55309 40885 55321 40888
rect 55355 40885 55367 40919
rect 55309 40879 55367 40885
rect 55674 40876 55680 40928
rect 55732 40876 55738 40928
rect 55766 40876 55772 40928
rect 55824 40876 55830 40928
rect 56134 40876 56140 40928
rect 56192 40876 56198 40928
rect 56336 40916 56364 40956
rect 56594 40944 56600 40996
rect 56652 40944 56658 40996
rect 57054 40944 57060 40996
rect 57112 40944 57118 40996
rect 57146 40916 57152 40928
rect 56336 40888 57152 40916
rect 57146 40876 57152 40888
rect 57204 40876 57210 40928
rect 57256 40916 57284 41024
rect 57606 41012 57612 41064
rect 57664 41012 57670 41064
rect 57793 41055 57851 41061
rect 57793 41021 57805 41055
rect 57839 41021 57851 41055
rect 60706 41052 60734 41160
rect 66070 41052 66076 41064
rect 60706 41024 66076 41052
rect 57793 41015 57851 41021
rect 57514 40944 57520 40996
rect 57572 40984 57578 40996
rect 57808 40984 57836 41015
rect 66070 41012 66076 41024
rect 66128 41012 66134 41064
rect 57572 40956 57836 40984
rect 57572 40944 57578 40956
rect 64874 40916 64880 40928
rect 57256 40888 64880 40916
rect 64874 40876 64880 40888
rect 64932 40876 64938 40928
rect 552 40826 66424 40848
rect 552 40774 2918 40826
rect 2970 40774 2982 40826
rect 3034 40774 3046 40826
rect 3098 40774 3110 40826
rect 3162 40774 3174 40826
rect 3226 40774 51918 40826
rect 51970 40774 51982 40826
rect 52034 40774 52046 40826
rect 52098 40774 52110 40826
rect 52162 40774 52174 40826
rect 52226 40774 66424 40826
rect 552 40752 66424 40774
rect 10686 40672 10692 40724
rect 10744 40712 10750 40724
rect 10965 40715 11023 40721
rect 10965 40712 10977 40715
rect 10744 40684 10977 40712
rect 10744 40672 10750 40684
rect 10965 40681 10977 40684
rect 11011 40681 11023 40715
rect 10965 40675 11023 40681
rect 11333 40715 11391 40721
rect 11333 40681 11345 40715
rect 11379 40712 11391 40715
rect 11422 40712 11428 40724
rect 11379 40684 11428 40712
rect 11379 40681 11391 40684
rect 11333 40675 11391 40681
rect 11422 40672 11428 40684
rect 11480 40672 11486 40724
rect 15933 40715 15991 40721
rect 15933 40681 15945 40715
rect 15979 40712 15991 40715
rect 16942 40712 16948 40724
rect 15979 40684 16948 40712
rect 15979 40681 15991 40684
rect 15933 40675 15991 40681
rect 16942 40672 16948 40684
rect 17000 40672 17006 40724
rect 17313 40715 17371 40721
rect 17313 40681 17325 40715
rect 17359 40712 17371 40715
rect 17865 40715 17923 40721
rect 17865 40712 17877 40715
rect 17359 40684 17877 40712
rect 17359 40681 17371 40684
rect 17313 40675 17371 40681
rect 17865 40681 17877 40684
rect 17911 40681 17923 40715
rect 20806 40712 20812 40724
rect 17865 40675 17923 40681
rect 19076 40684 20812 40712
rect 11532 40616 12926 40644
rect 10134 40536 10140 40588
rect 10192 40536 10198 40588
rect 10318 40536 10324 40588
rect 10376 40576 10382 40588
rect 10781 40579 10839 40585
rect 10781 40576 10793 40579
rect 10376 40548 10793 40576
rect 10376 40536 10382 40548
rect 10781 40545 10793 40548
rect 10827 40576 10839 40579
rect 11422 40576 11428 40588
rect 10827 40548 11428 40576
rect 10827 40545 10839 40548
rect 10781 40539 10839 40545
rect 11422 40536 11428 40548
rect 11480 40536 11486 40588
rect 8754 40468 8760 40520
rect 8812 40468 8818 40520
rect 9030 40468 9036 40520
rect 9088 40468 9094 40520
rect 9766 40468 9772 40520
rect 9824 40508 9830 40520
rect 10152 40508 10180 40536
rect 11532 40508 11560 40616
rect 14090 40604 14096 40656
rect 14148 40604 14154 40656
rect 15473 40647 15531 40653
rect 15473 40613 15485 40647
rect 15519 40644 15531 40647
rect 16758 40644 16764 40656
rect 15519 40616 16764 40644
rect 15519 40613 15531 40616
rect 15473 40607 15531 40613
rect 14369 40579 14427 40585
rect 14369 40545 14381 40579
rect 14415 40576 14427 40579
rect 15194 40576 15200 40588
rect 14415 40548 15200 40576
rect 14415 40545 14427 40548
rect 14369 40539 14427 40545
rect 15194 40536 15200 40548
rect 15252 40536 15258 40588
rect 9824 40480 11560 40508
rect 11609 40511 11667 40517
rect 9824 40468 9830 40480
rect 11609 40477 11621 40511
rect 11655 40508 11667 40511
rect 12250 40508 12256 40520
rect 11655 40480 12256 40508
rect 11655 40477 11667 40480
rect 11609 40471 11667 40477
rect 12250 40468 12256 40480
rect 12308 40468 12314 40520
rect 12345 40511 12403 40517
rect 12345 40477 12357 40511
rect 12391 40508 12403 40511
rect 13722 40508 13728 40520
rect 12391 40480 13728 40508
rect 12391 40477 12403 40480
rect 12345 40471 12403 40477
rect 13722 40468 13728 40480
rect 13780 40468 13786 40520
rect 14553 40511 14611 40517
rect 14553 40477 14565 40511
rect 14599 40477 14611 40511
rect 14553 40471 14611 40477
rect 14568 40440 14596 40471
rect 15378 40468 15384 40520
rect 15436 40468 15442 40520
rect 15488 40440 15516 40607
rect 16758 40604 16764 40616
rect 16816 40604 16822 40656
rect 17221 40647 17279 40653
rect 17221 40613 17233 40647
rect 17267 40644 17279 40647
rect 17402 40644 17408 40656
rect 17267 40616 17408 40644
rect 17267 40613 17279 40616
rect 17221 40607 17279 40613
rect 17402 40604 17408 40616
rect 17460 40604 17466 40656
rect 15565 40579 15623 40585
rect 15565 40545 15577 40579
rect 15611 40576 15623 40579
rect 17954 40576 17960 40588
rect 15611 40548 17960 40576
rect 15611 40545 15623 40548
rect 15565 40539 15623 40545
rect 17954 40536 17960 40548
rect 18012 40536 18018 40588
rect 19076 40585 19104 40684
rect 20806 40672 20812 40684
rect 20864 40672 20870 40724
rect 21266 40672 21272 40724
rect 21324 40672 21330 40724
rect 22186 40672 22192 40724
rect 22244 40672 22250 40724
rect 24762 40672 24768 40724
rect 24820 40712 24826 40724
rect 25501 40715 25559 40721
rect 25501 40712 25513 40715
rect 24820 40684 25513 40712
rect 24820 40672 24826 40684
rect 25501 40681 25513 40684
rect 25547 40681 25559 40715
rect 25501 40675 25559 40681
rect 26234 40672 26240 40724
rect 26292 40712 26298 40724
rect 26789 40715 26847 40721
rect 26789 40712 26801 40715
rect 26292 40684 26801 40712
rect 26292 40672 26298 40684
rect 26789 40681 26801 40684
rect 26835 40712 26847 40715
rect 26835 40684 27844 40712
rect 26835 40681 26847 40684
rect 26789 40675 26847 40681
rect 23934 40604 23940 40656
rect 23992 40604 23998 40656
rect 25222 40644 25228 40656
rect 25162 40616 25228 40644
rect 25222 40604 25228 40616
rect 25280 40604 25286 40656
rect 25869 40647 25927 40653
rect 25869 40613 25881 40647
rect 25915 40644 25927 40647
rect 27249 40647 27307 40653
rect 27249 40644 27261 40647
rect 25915 40616 27261 40644
rect 25915 40613 25927 40616
rect 25869 40607 25927 40613
rect 27249 40613 27261 40616
rect 27295 40613 27307 40647
rect 27249 40607 27307 40613
rect 18233 40579 18291 40585
rect 18233 40545 18245 40579
rect 18279 40545 18291 40579
rect 18233 40539 18291 40545
rect 19061 40579 19119 40585
rect 19061 40545 19073 40579
rect 19107 40545 19119 40579
rect 19061 40539 19119 40545
rect 16758 40468 16764 40520
rect 16816 40508 16822 40520
rect 17405 40511 17463 40517
rect 17405 40508 17417 40511
rect 16816 40480 17417 40508
rect 16816 40468 16822 40480
rect 17405 40477 17417 40480
rect 17451 40508 17463 40511
rect 17494 40508 17500 40520
rect 17451 40480 17500 40508
rect 17451 40477 17463 40480
rect 17405 40471 17463 40477
rect 17494 40468 17500 40480
rect 17552 40468 17558 40520
rect 17773 40511 17831 40517
rect 17773 40477 17785 40511
rect 17819 40508 17831 40511
rect 18046 40508 18052 40520
rect 17819 40480 18052 40508
rect 17819 40477 17831 40480
rect 17773 40471 17831 40477
rect 18046 40468 18052 40480
rect 18104 40508 18110 40520
rect 18248 40508 18276 40539
rect 20438 40536 20444 40588
rect 20496 40536 20502 40588
rect 21637 40579 21695 40585
rect 21637 40545 21649 40579
rect 21683 40576 21695 40579
rect 22830 40576 22836 40588
rect 21683 40548 22836 40576
rect 21683 40545 21695 40548
rect 21637 40539 21695 40545
rect 22830 40536 22836 40548
rect 22888 40536 22894 40588
rect 25961 40579 26019 40585
rect 25961 40545 25973 40579
rect 26007 40576 26019 40579
rect 26418 40576 26424 40588
rect 26007 40548 26424 40576
rect 26007 40545 26019 40548
rect 25961 40539 26019 40545
rect 26418 40536 26424 40548
rect 26476 40536 26482 40588
rect 26510 40536 26516 40588
rect 26568 40576 26574 40588
rect 27816 40585 27844 40684
rect 29086 40672 29092 40724
rect 29144 40672 29150 40724
rect 30558 40712 30564 40724
rect 30300 40684 30564 40712
rect 29914 40604 29920 40656
rect 29972 40604 29978 40656
rect 30006 40604 30012 40656
rect 30064 40644 30070 40656
rect 30300 40644 30328 40684
rect 30558 40672 30564 40684
rect 30616 40672 30622 40724
rect 30650 40672 30656 40724
rect 30708 40712 30714 40724
rect 31389 40715 31447 40721
rect 31389 40712 31401 40715
rect 30708 40684 31401 40712
rect 30708 40672 30714 40684
rect 31389 40681 31401 40684
rect 31435 40712 31447 40715
rect 32493 40715 32551 40721
rect 32493 40712 32505 40715
rect 31435 40684 32505 40712
rect 31435 40681 31447 40684
rect 31389 40675 31447 40681
rect 32493 40681 32505 40684
rect 32539 40681 32551 40715
rect 32493 40675 32551 40681
rect 32953 40715 33011 40721
rect 32953 40681 32965 40715
rect 32999 40712 33011 40715
rect 33226 40712 33232 40724
rect 32999 40684 33232 40712
rect 32999 40681 33011 40684
rect 32953 40675 33011 40681
rect 33226 40672 33232 40684
rect 33284 40672 33290 40724
rect 33686 40672 33692 40724
rect 33744 40712 33750 40724
rect 34149 40715 34207 40721
rect 34149 40712 34161 40715
rect 33744 40684 34161 40712
rect 33744 40672 33750 40684
rect 34149 40681 34161 40684
rect 34195 40681 34207 40715
rect 34149 40675 34207 40681
rect 34517 40715 34575 40721
rect 34517 40681 34529 40715
rect 34563 40712 34575 40715
rect 34606 40712 34612 40724
rect 34563 40684 34612 40712
rect 34563 40681 34575 40684
rect 34517 40675 34575 40681
rect 34606 40672 34612 40684
rect 34664 40672 34670 40724
rect 35894 40712 35900 40724
rect 34808 40684 35900 40712
rect 30064 40616 30406 40644
rect 30064 40604 30070 40616
rect 32122 40604 32128 40656
rect 32180 40644 32186 40656
rect 33042 40644 33048 40656
rect 32180 40616 33048 40644
rect 32180 40604 32186 40616
rect 33042 40604 33048 40616
rect 33100 40644 33106 40656
rect 34808 40644 34836 40684
rect 35894 40672 35900 40684
rect 35952 40672 35958 40724
rect 36538 40672 36544 40724
rect 36596 40672 36602 40724
rect 38562 40672 38568 40724
rect 38620 40712 38626 40724
rect 51166 40712 51172 40724
rect 38620 40684 51172 40712
rect 38620 40672 38626 40684
rect 33100 40616 34836 40644
rect 33100 40604 33106 40616
rect 27801 40579 27859 40585
rect 26568 40548 27568 40576
rect 26568 40536 26574 40548
rect 27540 40520 27568 40548
rect 27801 40545 27813 40579
rect 27847 40545 27859 40579
rect 27801 40539 27859 40545
rect 28721 40579 28779 40585
rect 28721 40545 28733 40579
rect 28767 40576 28779 40579
rect 28810 40576 28816 40588
rect 28767 40548 28816 40576
rect 28767 40545 28779 40548
rect 28721 40539 28779 40545
rect 28810 40536 28816 40548
rect 28868 40576 28874 40588
rect 29181 40579 29239 40585
rect 29181 40576 29193 40579
rect 28868 40548 29193 40576
rect 28868 40536 28874 40548
rect 29181 40545 29193 40548
rect 29227 40545 29239 40579
rect 29181 40539 29239 40545
rect 31662 40536 31668 40588
rect 31720 40536 31726 40588
rect 32585 40579 32643 40585
rect 32585 40545 32597 40579
rect 32631 40576 32643 40579
rect 33134 40576 33140 40588
rect 32631 40548 33140 40576
rect 32631 40545 32643 40548
rect 32585 40539 32643 40545
rect 33134 40536 33140 40548
rect 33192 40536 33198 40588
rect 33321 40579 33379 40585
rect 33321 40545 33333 40579
rect 33367 40545 33379 40579
rect 33321 40539 33379 40545
rect 33413 40579 33471 40585
rect 33413 40545 33425 40579
rect 33459 40576 33471 40579
rect 33778 40576 33784 40588
rect 33459 40548 33784 40576
rect 33459 40545 33471 40548
rect 33413 40539 33471 40545
rect 18104 40480 18276 40508
rect 18104 40468 18110 40480
rect 18322 40468 18328 40520
rect 18380 40468 18386 40520
rect 18414 40468 18420 40520
rect 18472 40468 18478 40520
rect 19334 40468 19340 40520
rect 19392 40468 19398 40520
rect 19886 40468 19892 40520
rect 19944 40508 19950 40520
rect 20346 40508 20352 40520
rect 19944 40480 20352 40508
rect 19944 40468 19950 40480
rect 20346 40468 20352 40480
rect 20404 40468 20410 40520
rect 20714 40468 20720 40520
rect 20772 40508 20778 40520
rect 21450 40508 21456 40520
rect 20772 40480 21456 40508
rect 20772 40468 20778 40480
rect 21450 40468 21456 40480
rect 21508 40468 21514 40520
rect 21729 40511 21787 40517
rect 21729 40477 21741 40511
rect 21775 40477 21787 40511
rect 21729 40471 21787 40477
rect 21913 40511 21971 40517
rect 21913 40477 21925 40511
rect 21959 40508 21971 40511
rect 22186 40508 22192 40520
rect 21959 40480 22192 40508
rect 21959 40477 21971 40480
rect 21913 40471 21971 40477
rect 21634 40440 21640 40452
rect 14568 40412 15516 40440
rect 20364 40412 21640 40440
rect 15105 40375 15163 40381
rect 15105 40341 15117 40375
rect 15151 40372 15163 40375
rect 15562 40372 15568 40384
rect 15151 40344 15568 40372
rect 15151 40341 15163 40344
rect 15105 40335 15163 40341
rect 15562 40332 15568 40344
rect 15620 40332 15626 40384
rect 16850 40332 16856 40384
rect 16908 40332 16914 40384
rect 17770 40332 17776 40384
rect 17828 40372 17834 40384
rect 20364 40372 20392 40412
rect 21634 40400 21640 40412
rect 21692 40400 21698 40452
rect 17828 40344 20392 40372
rect 17828 40332 17834 40344
rect 20622 40332 20628 40384
rect 20680 40372 20686 40384
rect 20809 40375 20867 40381
rect 20809 40372 20821 40375
rect 20680 40344 20821 40372
rect 20680 40332 20686 40344
rect 20809 40341 20821 40344
rect 20855 40372 20867 40375
rect 21744 40372 21772 40471
rect 22186 40468 22192 40480
rect 22244 40468 22250 40520
rect 23566 40468 23572 40520
rect 23624 40468 23630 40520
rect 23658 40468 23664 40520
rect 23716 40468 23722 40520
rect 25130 40508 25136 40520
rect 23768 40480 25136 40508
rect 23768 40440 23796 40480
rect 25130 40468 25136 40480
rect 25188 40468 25194 40520
rect 26053 40511 26111 40517
rect 26053 40508 26065 40511
rect 25332 40480 26065 40508
rect 22112 40412 23796 40440
rect 22112 40384 22140 40412
rect 20855 40344 21772 40372
rect 20855 40341 20867 40344
rect 20809 40335 20867 40341
rect 22094 40332 22100 40384
rect 22152 40332 22158 40384
rect 22922 40332 22928 40384
rect 22980 40332 22986 40384
rect 23290 40332 23296 40384
rect 23348 40372 23354 40384
rect 25332 40372 25360 40480
rect 26053 40477 26065 40480
rect 26099 40508 26111 40511
rect 26326 40508 26332 40520
rect 26099 40480 26332 40508
rect 26099 40477 26111 40480
rect 26053 40471 26111 40477
rect 26326 40468 26332 40480
rect 26384 40508 26390 40520
rect 26786 40508 26792 40520
rect 26384 40480 26792 40508
rect 26384 40468 26390 40480
rect 26786 40468 26792 40480
rect 26844 40468 26850 40520
rect 26878 40468 26884 40520
rect 26936 40468 26942 40520
rect 27062 40468 27068 40520
rect 27120 40468 27126 40520
rect 27522 40468 27528 40520
rect 27580 40508 27586 40520
rect 28997 40511 29055 40517
rect 28997 40508 29009 40511
rect 27580 40480 29009 40508
rect 27580 40468 27586 40480
rect 28997 40477 29009 40480
rect 29043 40508 29055 40511
rect 29270 40508 29276 40520
rect 29043 40480 29276 40508
rect 29043 40477 29055 40480
rect 28997 40471 29055 40477
rect 29270 40468 29276 40480
rect 29328 40468 29334 40520
rect 29362 40468 29368 40520
rect 29420 40508 29426 40520
rect 29641 40511 29699 40517
rect 29641 40508 29653 40511
rect 29420 40480 29653 40508
rect 29420 40468 29426 40480
rect 29641 40477 29653 40480
rect 29687 40477 29699 40511
rect 29641 40471 29699 40477
rect 30374 40468 30380 40520
rect 30432 40508 30438 40520
rect 30432 40480 30972 40508
rect 30432 40468 30438 40480
rect 26142 40400 26148 40452
rect 26200 40440 26206 40452
rect 30944 40440 30972 40480
rect 31202 40468 31208 40520
rect 31260 40508 31266 40520
rect 31846 40508 31852 40520
rect 31260 40480 31852 40508
rect 31260 40468 31266 40480
rect 31846 40468 31852 40480
rect 31904 40508 31910 40520
rect 32677 40511 32735 40517
rect 32677 40508 32689 40511
rect 31904 40480 32689 40508
rect 31904 40468 31910 40480
rect 32677 40477 32689 40480
rect 32723 40477 32735 40511
rect 32677 40471 32735 40477
rect 32950 40468 32956 40520
rect 33008 40508 33014 40520
rect 33336 40508 33364 40539
rect 33778 40536 33784 40548
rect 33836 40536 33842 40588
rect 34808 40585 34836 40616
rect 35066 40604 35072 40656
rect 35124 40604 35130 40656
rect 35526 40604 35532 40656
rect 35584 40604 35590 40656
rect 37550 40604 37556 40656
rect 37608 40644 37614 40656
rect 37645 40647 37703 40653
rect 37645 40644 37657 40647
rect 37608 40616 37657 40644
rect 37608 40604 37614 40616
rect 37645 40613 37657 40616
rect 37691 40613 37703 40647
rect 39022 40644 39028 40656
rect 38870 40616 39028 40644
rect 37645 40607 37703 40613
rect 39022 40604 39028 40616
rect 39080 40604 39086 40656
rect 40034 40644 40040 40656
rect 39500 40616 40040 40644
rect 34793 40579 34851 40585
rect 34793 40545 34805 40579
rect 34839 40545 34851 40579
rect 34793 40539 34851 40545
rect 37182 40536 37188 40588
rect 37240 40576 37246 40588
rect 37369 40579 37427 40585
rect 37369 40576 37381 40579
rect 37240 40548 37381 40576
rect 37240 40536 37246 40548
rect 37369 40545 37381 40548
rect 37415 40545 37427 40579
rect 39500 40576 39528 40616
rect 40034 40604 40040 40616
rect 40092 40604 40098 40656
rect 40770 40604 40776 40656
rect 40828 40644 40834 40656
rect 41322 40644 41328 40656
rect 40828 40616 41328 40644
rect 40828 40604 40834 40616
rect 41322 40604 41328 40616
rect 41380 40604 41386 40656
rect 41892 40653 41920 40684
rect 51166 40672 51172 40684
rect 51224 40672 51230 40724
rect 51261 40715 51319 40721
rect 51261 40681 51273 40715
rect 51307 40712 51319 40715
rect 51442 40712 51448 40724
rect 51307 40684 51448 40712
rect 51307 40681 51319 40684
rect 51261 40675 51319 40681
rect 51442 40672 51448 40684
rect 51500 40672 51506 40724
rect 52362 40672 52368 40724
rect 52420 40712 52426 40724
rect 52420 40684 54892 40712
rect 52420 40672 52426 40684
rect 41877 40647 41935 40653
rect 41877 40613 41889 40647
rect 41923 40613 41935 40647
rect 41877 40607 41935 40613
rect 44726 40604 44732 40656
rect 44784 40644 44790 40656
rect 44784 40616 45600 40644
rect 44784 40604 44790 40616
rect 37369 40539 37427 40545
rect 39132 40548 39528 40576
rect 39577 40579 39635 40585
rect 33008 40480 33364 40508
rect 33008 40468 33014 40480
rect 33502 40468 33508 40520
rect 33560 40508 33566 40520
rect 33597 40511 33655 40517
rect 33597 40508 33609 40511
rect 33560 40480 33609 40508
rect 33560 40468 33566 40480
rect 33597 40477 33609 40480
rect 33643 40508 33655 40511
rect 33962 40508 33968 40520
rect 33643 40480 33968 40508
rect 33643 40477 33655 40480
rect 33597 40471 33655 40477
rect 33962 40468 33968 40480
rect 34020 40468 34026 40520
rect 34054 40468 34060 40520
rect 34112 40468 34118 40520
rect 36078 40468 36084 40520
rect 36136 40508 36142 40520
rect 37642 40508 37648 40520
rect 36136 40480 37648 40508
rect 36136 40468 36142 40480
rect 37642 40468 37648 40480
rect 37700 40468 37706 40520
rect 38378 40468 38384 40520
rect 38436 40508 38442 40520
rect 39132 40517 39160 40548
rect 39577 40545 39589 40579
rect 39623 40576 39635 40579
rect 40126 40576 40132 40588
rect 39623 40548 40132 40576
rect 39623 40545 39635 40548
rect 39577 40539 39635 40545
rect 40126 40536 40132 40548
rect 40184 40536 40190 40588
rect 40681 40579 40739 40585
rect 40681 40545 40693 40579
rect 40727 40576 40739 40579
rect 40954 40576 40960 40588
rect 40727 40548 40960 40576
rect 40727 40545 40739 40548
rect 40681 40539 40739 40545
rect 40954 40536 40960 40548
rect 41012 40536 41018 40588
rect 41601 40579 41659 40585
rect 41601 40545 41613 40579
rect 41647 40576 41659 40579
rect 41966 40576 41972 40588
rect 41647 40548 41972 40576
rect 41647 40545 41659 40548
rect 41601 40539 41659 40545
rect 39117 40511 39175 40517
rect 38436 40480 38700 40508
rect 38436 40468 38442 40480
rect 38672 40440 38700 40480
rect 39117 40477 39129 40511
rect 39163 40477 39175 40511
rect 39117 40471 39175 40477
rect 39298 40468 39304 40520
rect 39356 40508 39362 40520
rect 39669 40511 39727 40517
rect 39669 40508 39681 40511
rect 39356 40480 39681 40508
rect 39356 40468 39362 40480
rect 39669 40477 39681 40480
rect 39715 40477 39727 40511
rect 39669 40471 39727 40477
rect 39761 40511 39819 40517
rect 39761 40477 39773 40511
rect 39807 40477 39819 40511
rect 39761 40471 39819 40477
rect 39776 40440 39804 40471
rect 39850 40468 39856 40520
rect 39908 40508 39914 40520
rect 40773 40511 40831 40517
rect 40773 40508 40785 40511
rect 39908 40480 40785 40508
rect 39908 40468 39914 40480
rect 40773 40477 40785 40480
rect 40819 40477 40831 40511
rect 40773 40471 40831 40477
rect 40865 40511 40923 40517
rect 40865 40477 40877 40511
rect 40911 40477 40923 40511
rect 40865 40471 40923 40477
rect 26200 40412 29684 40440
rect 30944 40412 34928 40440
rect 38672 40412 39804 40440
rect 26200 40400 26206 40412
rect 23348 40344 25360 40372
rect 25409 40375 25467 40381
rect 23348 40332 23354 40344
rect 25409 40341 25421 40375
rect 25455 40372 25467 40375
rect 25590 40372 25596 40384
rect 25455 40344 25596 40372
rect 25455 40341 25467 40344
rect 25409 40335 25467 40341
rect 25590 40332 25596 40344
rect 25648 40332 25654 40384
rect 26421 40375 26479 40381
rect 26421 40341 26433 40375
rect 26467 40372 26479 40375
rect 26694 40372 26700 40384
rect 26467 40344 26700 40372
rect 26467 40341 26479 40344
rect 26421 40335 26479 40341
rect 26694 40332 26700 40344
rect 26752 40332 26758 40384
rect 28074 40332 28080 40384
rect 28132 40332 28138 40384
rect 29270 40332 29276 40384
rect 29328 40372 29334 40384
rect 29549 40375 29607 40381
rect 29549 40372 29561 40375
rect 29328 40344 29561 40372
rect 29328 40332 29334 40344
rect 29549 40341 29561 40344
rect 29595 40341 29607 40375
rect 29656 40372 29684 40412
rect 30466 40372 30472 40384
rect 29656 40344 30472 40372
rect 29549 40335 29607 40341
rect 30466 40332 30472 40344
rect 30524 40332 30530 40384
rect 31846 40332 31852 40384
rect 31904 40372 31910 40384
rect 31941 40375 31999 40381
rect 31941 40372 31953 40375
rect 31904 40344 31953 40372
rect 31904 40332 31910 40344
rect 31941 40341 31953 40344
rect 31987 40341 31999 40375
rect 31941 40335 31999 40341
rect 32122 40332 32128 40384
rect 32180 40332 32186 40384
rect 34900 40372 34928 40412
rect 40310 40400 40316 40452
rect 40368 40400 40374 40452
rect 40678 40400 40684 40452
rect 40736 40440 40742 40452
rect 40880 40440 40908 40471
rect 40736 40412 40908 40440
rect 40736 40400 40742 40412
rect 38654 40372 38660 40384
rect 34900 40344 38660 40372
rect 38654 40332 38660 40344
rect 38712 40332 38718 40384
rect 39206 40332 39212 40384
rect 39264 40332 39270 40384
rect 40402 40332 40408 40384
rect 40460 40372 40466 40384
rect 41616 40372 41644 40539
rect 41966 40536 41972 40548
rect 42024 40536 42030 40588
rect 45462 40536 45468 40588
rect 45520 40536 45526 40588
rect 45572 40576 45600 40616
rect 45738 40604 45744 40656
rect 45796 40644 45802 40656
rect 45925 40647 45983 40653
rect 45925 40644 45937 40647
rect 45796 40616 45937 40644
rect 45796 40604 45802 40616
rect 45925 40613 45937 40616
rect 45971 40613 45983 40647
rect 45925 40607 45983 40613
rect 46382 40604 46388 40656
rect 46440 40644 46446 40656
rect 47397 40647 47455 40653
rect 47397 40644 47409 40647
rect 46440 40616 47409 40644
rect 46440 40604 46446 40616
rect 47397 40613 47409 40616
rect 47443 40613 47455 40647
rect 47397 40607 47455 40613
rect 49418 40604 49424 40656
rect 49476 40604 49482 40656
rect 49970 40604 49976 40656
rect 50028 40604 50034 40656
rect 50706 40604 50712 40656
rect 50764 40644 50770 40656
rect 51629 40647 51687 40653
rect 51629 40644 51641 40647
rect 50764 40616 51641 40644
rect 50764 40604 50770 40616
rect 51629 40613 51641 40616
rect 51675 40613 51687 40647
rect 51629 40607 51687 40613
rect 51736 40616 53052 40644
rect 46198 40576 46204 40588
rect 45572 40548 46204 40576
rect 46198 40536 46204 40548
rect 46256 40536 46262 40588
rect 47489 40579 47547 40585
rect 47489 40545 47501 40579
rect 47535 40576 47547 40579
rect 47670 40576 47676 40588
rect 47535 40548 47676 40576
rect 47535 40545 47547 40548
rect 47489 40539 47547 40545
rect 47670 40536 47676 40548
rect 47728 40536 47734 40588
rect 47762 40536 47768 40588
rect 47820 40576 47826 40588
rect 48222 40576 48228 40588
rect 47820 40548 48228 40576
rect 47820 40536 47826 40548
rect 48222 40536 48228 40548
rect 48280 40536 48286 40588
rect 51074 40536 51080 40588
rect 51132 40576 51138 40588
rect 51736 40576 51764 40616
rect 51132 40548 51764 40576
rect 51132 40536 51138 40548
rect 52270 40536 52276 40588
rect 52328 40576 52334 40588
rect 52457 40579 52515 40585
rect 52457 40576 52469 40579
rect 52328 40548 52469 40576
rect 52328 40536 52334 40548
rect 52457 40545 52469 40548
rect 52503 40545 52515 40579
rect 52457 40539 52515 40545
rect 43714 40468 43720 40520
rect 43772 40468 43778 40520
rect 45189 40511 45247 40517
rect 45189 40477 45201 40511
rect 45235 40508 45247 40511
rect 46017 40511 46075 40517
rect 45235 40480 45600 40508
rect 45235 40477 45247 40480
rect 45189 40471 45247 40477
rect 45572 40449 45600 40480
rect 46017 40477 46029 40511
rect 46063 40477 46075 40511
rect 46017 40471 46075 40477
rect 46109 40511 46167 40517
rect 46109 40477 46121 40511
rect 46155 40508 46167 40511
rect 47581 40511 47639 40517
rect 46155 40480 47348 40508
rect 46155 40477 46167 40480
rect 46109 40471 46167 40477
rect 45557 40443 45615 40449
rect 45557 40409 45569 40443
rect 45603 40409 45615 40443
rect 46032 40440 46060 40471
rect 47029 40443 47087 40449
rect 47029 40440 47041 40443
rect 46032 40412 47041 40440
rect 45557 40403 45615 40409
rect 47029 40409 47041 40412
rect 47075 40409 47087 40443
rect 47029 40403 47087 40409
rect 40460 40344 41644 40372
rect 40460 40332 40466 40344
rect 43346 40332 43352 40384
rect 43404 40332 43410 40384
rect 47320 40372 47348 40480
rect 47581 40477 47593 40511
rect 47627 40508 47639 40511
rect 47854 40508 47860 40520
rect 47627 40480 47860 40508
rect 47627 40477 47639 40480
rect 47581 40471 47639 40477
rect 47854 40468 47860 40480
rect 47912 40468 47918 40520
rect 48498 40468 48504 40520
rect 48556 40468 48562 40520
rect 49145 40511 49203 40517
rect 49145 40477 49157 40511
rect 49191 40477 49203 40511
rect 49145 40471 49203 40477
rect 47394 40400 47400 40452
rect 47452 40440 47458 40452
rect 48222 40440 48228 40452
rect 47452 40412 48228 40440
rect 47452 40400 47458 40412
rect 48222 40400 48228 40412
rect 48280 40440 48286 40452
rect 49160 40440 49188 40471
rect 50154 40468 50160 40520
rect 50212 40508 50218 40520
rect 50706 40508 50712 40520
rect 50212 40480 50712 40508
rect 50212 40468 50218 40480
rect 50706 40468 50712 40480
rect 50764 40508 50770 40520
rect 51169 40511 51227 40517
rect 51169 40508 51181 40511
rect 50764 40480 51181 40508
rect 50764 40468 50770 40480
rect 51169 40477 51181 40480
rect 51215 40508 51227 40511
rect 51721 40511 51779 40517
rect 51721 40508 51733 40511
rect 51215 40480 51733 40508
rect 51215 40477 51227 40480
rect 51169 40471 51227 40477
rect 51721 40477 51733 40480
rect 51767 40477 51779 40511
rect 51721 40471 51779 40477
rect 51810 40468 51816 40520
rect 51868 40468 51874 40520
rect 52822 40468 52828 40520
rect 52880 40468 52886 40520
rect 53024 40508 53052 40616
rect 53466 40536 53472 40588
rect 53524 40536 53530 40588
rect 54864 40585 54892 40684
rect 55122 40672 55128 40724
rect 55180 40712 55186 40724
rect 55180 40684 55352 40712
rect 55180 40672 55186 40684
rect 55214 40604 55220 40656
rect 55272 40604 55278 40656
rect 55324 40644 55352 40684
rect 56686 40672 56692 40724
rect 56744 40712 56750 40724
rect 57514 40712 57520 40724
rect 56744 40684 57520 40712
rect 56744 40672 56750 40684
rect 57514 40672 57520 40684
rect 57572 40672 57578 40724
rect 57698 40672 57704 40724
rect 57756 40712 57762 40724
rect 60642 40712 60648 40724
rect 57756 40684 60648 40712
rect 57756 40672 57762 40684
rect 60642 40672 60648 40684
rect 60700 40672 60706 40724
rect 55324 40616 55706 40644
rect 54849 40579 54907 40585
rect 54849 40545 54861 40579
rect 54895 40576 54907 40579
rect 54941 40579 54999 40585
rect 54941 40576 54953 40579
rect 54895 40548 54953 40576
rect 54895 40545 54907 40548
rect 54849 40539 54907 40545
rect 54941 40545 54953 40548
rect 54987 40545 54999 40579
rect 54941 40539 54999 40545
rect 54202 40508 54208 40520
rect 53024 40480 54208 40508
rect 54202 40468 54208 40480
rect 54260 40468 54266 40520
rect 54570 40468 54576 40520
rect 54628 40468 54634 40520
rect 55766 40468 55772 40520
rect 55824 40508 55830 40520
rect 56965 40511 57023 40517
rect 56965 40508 56977 40511
rect 55824 40480 56977 40508
rect 55824 40468 55830 40480
rect 56965 40477 56977 40480
rect 57011 40477 57023 40511
rect 56965 40471 57023 40477
rect 51350 40440 51356 40452
rect 48280 40412 49188 40440
rect 48280 40400 48286 40412
rect 47762 40372 47768 40384
rect 47320 40344 47768 40372
rect 47762 40332 47768 40344
rect 47820 40332 47826 40384
rect 49050 40332 49056 40384
rect 49108 40332 49114 40384
rect 49160 40372 49188 40412
rect 51046 40412 51356 40440
rect 51046 40372 51074 40412
rect 51350 40400 51356 40412
rect 51408 40400 51414 40452
rect 49160 40344 51074 40372
rect 52641 40375 52699 40381
rect 52641 40341 52653 40375
rect 52687 40372 52699 40375
rect 53558 40372 53564 40384
rect 52687 40344 53564 40372
rect 52687 40341 52699 40344
rect 52641 40335 52699 40341
rect 53558 40332 53564 40344
rect 53616 40332 53622 40384
rect 54478 40332 54484 40384
rect 54536 40372 54542 40384
rect 56686 40372 56692 40384
rect 54536 40344 56692 40372
rect 54536 40332 54542 40344
rect 56686 40332 56692 40344
rect 56744 40332 56750 40384
rect 552 40282 66424 40304
rect 552 40230 1998 40282
rect 2050 40230 2062 40282
rect 2114 40230 2126 40282
rect 2178 40230 2190 40282
rect 2242 40230 2254 40282
rect 2306 40230 50998 40282
rect 51050 40230 51062 40282
rect 51114 40230 51126 40282
rect 51178 40230 51190 40282
rect 51242 40230 51254 40282
rect 51306 40230 66424 40282
rect 552 40208 66424 40230
rect 9030 40128 9036 40180
rect 9088 40168 9094 40180
rect 9493 40171 9551 40177
rect 9493 40168 9505 40171
rect 9088 40140 9505 40168
rect 9088 40128 9094 40140
rect 9493 40137 9505 40140
rect 9539 40137 9551 40171
rect 10962 40168 10968 40180
rect 9493 40131 9551 40137
rect 9876 40140 10968 40168
rect 9876 40100 9904 40140
rect 10318 40100 10324 40112
rect 9324 40072 9904 40100
rect 9968 40072 10324 40100
rect 9324 40044 9352 40072
rect 9306 39992 9312 40044
rect 9364 39992 9370 40044
rect 9968 40041 9996 40072
rect 10318 40060 10324 40072
rect 10376 40060 10382 40112
rect 9953 40035 10011 40041
rect 9953 40001 9965 40035
rect 9999 40001 10011 40035
rect 9953 39995 10011 40001
rect 10137 40035 10195 40041
rect 10137 40001 10149 40035
rect 10183 40032 10195 40035
rect 10410 40032 10416 40044
rect 10183 40004 10416 40032
rect 10183 40001 10195 40004
rect 10137 39995 10195 40001
rect 10410 39992 10416 40004
rect 10468 39992 10474 40044
rect 10888 40041 10916 40140
rect 10962 40128 10968 40140
rect 11020 40128 11026 40180
rect 16288 40171 16346 40177
rect 13372 40140 16160 40168
rect 13372 40100 13400 40140
rect 11808 40072 13400 40100
rect 11808 40041 11836 40072
rect 10873 40035 10931 40041
rect 10873 40001 10885 40035
rect 10919 40001 10931 40035
rect 10873 39995 10931 40001
rect 11793 40035 11851 40041
rect 11793 40001 11805 40035
rect 11839 40001 11851 40035
rect 11793 39995 11851 40001
rect 12802 39992 12808 40044
rect 12860 40032 12866 40044
rect 13280 40041 13308 40072
rect 13081 40035 13139 40041
rect 13081 40032 13093 40035
rect 12860 40004 13093 40032
rect 12860 39992 12866 40004
rect 13081 40001 13093 40004
rect 13127 40001 13139 40035
rect 13081 39995 13139 40001
rect 13265 40035 13323 40041
rect 13265 40001 13277 40035
rect 13311 40001 13323 40035
rect 13265 39995 13323 40001
rect 14182 39992 14188 40044
rect 14240 39992 14246 40044
rect 14458 39992 14464 40044
rect 14516 39992 14522 40044
rect 15194 39992 15200 40044
rect 15252 40032 15258 40044
rect 16025 40035 16083 40041
rect 16025 40032 16037 40035
rect 15252 40004 16037 40032
rect 15252 39992 15258 40004
rect 16025 40001 16037 40004
rect 16071 40001 16083 40035
rect 16132 40032 16160 40140
rect 16288 40137 16300 40171
rect 16334 40168 16346 40171
rect 16850 40168 16856 40180
rect 16334 40140 16856 40168
rect 16334 40137 16346 40140
rect 16288 40131 16346 40137
rect 16850 40128 16856 40140
rect 16908 40128 16914 40180
rect 19794 40128 19800 40180
rect 19852 40168 19858 40180
rect 20438 40168 20444 40180
rect 19852 40140 20444 40168
rect 19852 40128 19858 40140
rect 20438 40128 20444 40140
rect 20496 40128 20502 40180
rect 20551 40171 20609 40177
rect 20551 40137 20563 40171
rect 20597 40168 20609 40171
rect 20901 40171 20959 40177
rect 20901 40168 20913 40171
rect 20597 40140 20913 40168
rect 20597 40137 20609 40140
rect 20551 40131 20609 40137
rect 20901 40137 20913 40140
rect 20947 40137 20959 40171
rect 20901 40131 20959 40137
rect 22097 40171 22155 40177
rect 22097 40137 22109 40171
rect 22143 40168 22155 40171
rect 22278 40168 22284 40180
rect 22143 40140 22284 40168
rect 22143 40137 22155 40140
rect 22097 40131 22155 40137
rect 22278 40128 22284 40140
rect 22336 40128 22342 40180
rect 23934 40128 23940 40180
rect 23992 40168 23998 40180
rect 24121 40171 24179 40177
rect 24121 40168 24133 40171
rect 23992 40140 24133 40168
rect 23992 40128 23998 40140
rect 24121 40137 24133 40140
rect 24167 40137 24179 40171
rect 26510 40168 26516 40180
rect 24121 40131 24179 40137
rect 24780 40140 26516 40168
rect 21082 40060 21088 40112
rect 21140 40100 21146 40112
rect 21140 40072 21496 40100
rect 21140 40060 21146 40072
rect 17310 40032 17316 40044
rect 16132 40004 17316 40032
rect 16025 39995 16083 40001
rect 17310 39992 17316 40004
rect 17368 39992 17374 40044
rect 17773 40035 17831 40041
rect 17773 40001 17785 40035
rect 17819 40032 17831 40035
rect 17954 40032 17960 40044
rect 17819 40004 17960 40032
rect 17819 40001 17831 40004
rect 17773 39995 17831 40001
rect 17954 39992 17960 40004
rect 18012 39992 18018 40044
rect 20070 39992 20076 40044
rect 20128 40032 20134 40044
rect 21468 40041 21496 40072
rect 21634 40060 21640 40112
rect 21692 40100 21698 40112
rect 21692 40072 22140 40100
rect 21692 40060 21698 40072
rect 22112 40044 22140 40072
rect 22186 40060 22192 40112
rect 22244 40100 22250 40112
rect 22244 40072 22692 40100
rect 22244 40060 22250 40072
rect 20809 40035 20867 40041
rect 20809 40032 20821 40035
rect 20128 40004 20821 40032
rect 20128 39992 20134 40004
rect 20809 40001 20821 40004
rect 20855 40001 20867 40035
rect 20809 39995 20867 40001
rect 21453 40035 21511 40041
rect 21453 40001 21465 40035
rect 21499 40001 21511 40035
rect 21453 39995 21511 40001
rect 22094 39992 22100 40044
rect 22152 39992 22158 40044
rect 22554 39992 22560 40044
rect 22612 39992 22618 40044
rect 22664 40041 22692 40072
rect 23290 40060 23296 40112
rect 23348 40100 23354 40112
rect 23348 40072 23520 40100
rect 23348 40060 23354 40072
rect 23492 40041 23520 40072
rect 24486 40060 24492 40112
rect 24544 40100 24550 40112
rect 24780 40100 24808 40140
rect 26510 40128 26516 40140
rect 26568 40128 26574 40180
rect 26694 40128 26700 40180
rect 26752 40177 26758 40180
rect 26752 40171 26767 40177
rect 26755 40137 26767 40171
rect 27982 40168 27988 40180
rect 26752 40131 26767 40137
rect 26896 40140 27988 40168
rect 26752 40128 26758 40131
rect 24544 40072 24808 40100
rect 24544 40060 24550 40072
rect 22649 40035 22707 40041
rect 22649 40001 22661 40035
rect 22695 40001 22707 40035
rect 22649 39995 22707 40001
rect 23477 40035 23535 40041
rect 23477 40001 23489 40035
rect 23523 40001 23535 40035
rect 23477 39995 23535 40001
rect 24394 39992 24400 40044
rect 24452 40032 24458 40044
rect 24780 40041 24808 40072
rect 24581 40035 24639 40041
rect 24581 40032 24593 40035
rect 24452 40004 24593 40032
rect 24452 39992 24458 40004
rect 24581 40001 24593 40004
rect 24627 40001 24639 40035
rect 24581 39995 24639 40001
rect 24765 40035 24823 40041
rect 24765 40001 24777 40035
rect 24811 40001 24823 40035
rect 26896 40032 26924 40140
rect 27982 40128 27988 40140
rect 28040 40128 28046 40180
rect 28810 40128 28816 40180
rect 28868 40128 28874 40180
rect 30282 40168 30288 40180
rect 29748 40140 30288 40168
rect 26970 40060 26976 40112
rect 27028 40060 27034 40112
rect 29748 40100 29776 40140
rect 30282 40128 30288 40140
rect 30340 40128 30346 40180
rect 30466 40128 30472 40180
rect 30524 40168 30530 40180
rect 36078 40168 36084 40180
rect 30524 40140 36084 40168
rect 30524 40128 30530 40140
rect 36078 40128 36084 40140
rect 36136 40128 36142 40180
rect 36262 40128 36268 40180
rect 36320 40168 36326 40180
rect 36722 40168 36728 40180
rect 36320 40140 36728 40168
rect 36320 40128 36326 40140
rect 36722 40128 36728 40140
rect 36780 40168 36786 40180
rect 37632 40171 37690 40177
rect 36780 40140 37228 40168
rect 36780 40128 36786 40140
rect 29656 40072 29776 40100
rect 24765 39995 24823 40001
rect 25608 40004 26924 40032
rect 26988 40032 27016 40060
rect 27065 40035 27123 40041
rect 27065 40032 27077 40035
rect 26988 40004 27077 40032
rect 7926 39924 7932 39976
rect 7984 39964 7990 39976
rect 12434 39964 12440 39976
rect 7984 39936 12440 39964
rect 7984 39924 7990 39936
rect 12434 39924 12440 39936
rect 12492 39924 12498 39976
rect 12989 39967 13047 39973
rect 12989 39933 13001 39967
rect 13035 39964 13047 39967
rect 13722 39964 13728 39976
rect 13035 39936 13728 39964
rect 13035 39933 13047 39936
rect 12989 39927 13047 39933
rect 13722 39924 13728 39936
rect 13780 39924 13786 39976
rect 20990 39924 20996 39976
rect 21048 39964 21054 39976
rect 21269 39967 21327 39973
rect 21269 39964 21281 39967
rect 21048 39936 21281 39964
rect 21048 39924 21054 39936
rect 21269 39933 21281 39936
rect 21315 39933 21327 39967
rect 21269 39927 21327 39933
rect 22922 39924 22928 39976
rect 22980 39964 22986 39976
rect 23293 39967 23351 39973
rect 23293 39964 23305 39967
rect 22980 39936 23305 39964
rect 22980 39924 22986 39936
rect 23293 39933 23305 39936
rect 23339 39933 23351 39967
rect 23293 39927 23351 39933
rect 23566 39924 23572 39976
rect 23624 39964 23630 39976
rect 24210 39964 24216 39976
rect 23624 39936 24216 39964
rect 23624 39924 23630 39936
rect 24210 39924 24216 39936
rect 24268 39964 24274 39976
rect 24489 39967 24547 39973
rect 24489 39964 24501 39967
rect 24268 39936 24501 39964
rect 24268 39924 24274 39936
rect 24489 39933 24501 39936
rect 24535 39933 24547 39967
rect 24489 39927 24547 39933
rect 25406 39924 25412 39976
rect 25464 39964 25470 39976
rect 25608 39964 25636 40004
rect 27065 40001 27077 40004
rect 27111 40032 27123 40035
rect 29362 40032 29368 40044
rect 27111 40004 29368 40032
rect 27111 40001 27123 40004
rect 27065 39995 27123 40001
rect 29362 39992 29368 40004
rect 29420 39992 29426 40044
rect 29656 40041 29684 40072
rect 31570 40060 31576 40112
rect 31628 40100 31634 40112
rect 35250 40100 35256 40112
rect 31628 40072 35256 40100
rect 31628 40060 31634 40072
rect 35250 40060 35256 40072
rect 35308 40060 35314 40112
rect 37200 40100 37228 40140
rect 37632 40137 37644 40171
rect 37678 40168 37690 40171
rect 39206 40168 39212 40180
rect 37678 40140 39212 40168
rect 37678 40137 37690 40140
rect 37632 40131 37690 40137
rect 39206 40128 39212 40140
rect 39264 40128 39270 40180
rect 39390 40128 39396 40180
rect 39448 40168 39454 40180
rect 41598 40168 41604 40180
rect 39448 40140 41604 40168
rect 39448 40128 39454 40140
rect 41598 40128 41604 40140
rect 41656 40168 41662 40180
rect 41874 40168 41880 40180
rect 41656 40140 41880 40168
rect 41656 40128 41662 40140
rect 41874 40128 41880 40140
rect 41932 40128 41938 40180
rect 46290 40128 46296 40180
rect 46348 40168 46354 40180
rect 46673 40171 46731 40177
rect 46673 40168 46685 40171
rect 46348 40140 46685 40168
rect 46348 40128 46354 40140
rect 46673 40137 46685 40140
rect 46719 40137 46731 40171
rect 48038 40168 48044 40180
rect 46673 40131 46731 40137
rect 46860 40140 48044 40168
rect 37200 40072 37320 40100
rect 29641 40035 29699 40041
rect 29641 40001 29653 40035
rect 29687 40001 29699 40035
rect 29641 39995 29699 40001
rect 29825 40035 29883 40041
rect 29825 40001 29837 40035
rect 29871 40032 29883 40035
rect 30098 40032 30104 40044
rect 29871 40004 30104 40032
rect 29871 40001 29883 40004
rect 29825 39995 29883 40001
rect 30098 39992 30104 40004
rect 30156 39992 30162 40044
rect 30558 39992 30564 40044
rect 30616 40032 30622 40044
rect 31294 40032 31300 40044
rect 30616 40004 31300 40032
rect 30616 39992 30622 40004
rect 31294 39992 31300 40004
rect 31352 39992 31358 40044
rect 31386 39992 31392 40044
rect 31444 40032 31450 40044
rect 36446 40032 36452 40044
rect 31444 40004 36452 40032
rect 31444 39992 31450 40004
rect 36446 39992 36452 40004
rect 36504 39992 36510 40044
rect 37093 40035 37151 40041
rect 37093 40001 37105 40035
rect 37139 40032 37151 40035
rect 37182 40032 37188 40044
rect 37139 40004 37188 40032
rect 37139 40001 37151 40004
rect 37093 39995 37151 40001
rect 37182 39992 37188 40004
rect 37240 39992 37246 40044
rect 37292 40032 37320 40072
rect 39040 40072 39528 40100
rect 37369 40035 37427 40041
rect 37369 40032 37381 40035
rect 37292 40004 37381 40032
rect 37369 40001 37381 40004
rect 37415 40001 37427 40035
rect 37369 39995 37427 40001
rect 38286 39992 38292 40044
rect 38344 40032 38350 40044
rect 39040 40032 39068 40072
rect 39500 40044 39528 40072
rect 44192 40072 45692 40100
rect 38344 40004 39068 40032
rect 39117 40035 39175 40041
rect 38344 39992 38350 40004
rect 39117 40001 39129 40035
rect 39163 40001 39175 40035
rect 39117 39995 39175 40001
rect 25464 39950 25636 39964
rect 26973 39967 27031 39973
rect 25464 39936 25622 39950
rect 25464 39924 25470 39936
rect 26973 39933 26985 39967
rect 27019 39933 27031 39967
rect 39022 39964 39028 39976
rect 38778 39936 39028 39964
rect 26973 39927 27031 39933
rect 8938 39856 8944 39908
rect 8996 39896 9002 39908
rect 9033 39899 9091 39905
rect 9033 39896 9045 39899
rect 8996 39868 9045 39896
rect 8996 39856 9002 39868
rect 9033 39865 9045 39868
rect 9079 39865 9091 39899
rect 9033 39859 9091 39865
rect 9125 39899 9183 39905
rect 9125 39865 9137 39899
rect 9171 39896 9183 39899
rect 9171 39868 11192 39896
rect 9171 39865 9183 39868
rect 9125 39859 9183 39865
rect 8202 39788 8208 39840
rect 8260 39828 8266 39840
rect 8665 39831 8723 39837
rect 8665 39828 8677 39831
rect 8260 39800 8677 39828
rect 8260 39788 8266 39800
rect 8665 39797 8677 39800
rect 8711 39797 8723 39831
rect 8665 39791 8723 39797
rect 9674 39788 9680 39840
rect 9732 39828 9738 39840
rect 9861 39831 9919 39837
rect 9861 39828 9873 39831
rect 9732 39800 9873 39828
rect 9732 39788 9738 39800
rect 9861 39797 9873 39800
rect 9907 39797 9919 39831
rect 9861 39791 9919 39797
rect 10134 39788 10140 39840
rect 10192 39828 10198 39840
rect 10321 39831 10379 39837
rect 10321 39828 10333 39831
rect 10192 39800 10333 39828
rect 10192 39788 10198 39800
rect 10321 39797 10333 39800
rect 10367 39797 10379 39831
rect 10321 39791 10379 39797
rect 10686 39788 10692 39840
rect 10744 39788 10750 39840
rect 10781 39831 10839 39837
rect 10781 39797 10793 39831
rect 10827 39828 10839 39831
rect 11054 39828 11060 39840
rect 10827 39800 11060 39828
rect 10827 39797 10839 39800
rect 10781 39791 10839 39797
rect 11054 39788 11060 39800
rect 11112 39788 11118 39840
rect 11164 39837 11192 39868
rect 11422 39856 11428 39908
rect 11480 39896 11486 39908
rect 11517 39899 11575 39905
rect 11517 39896 11529 39899
rect 11480 39868 11529 39896
rect 11480 39856 11486 39868
rect 11517 39865 11529 39868
rect 11563 39865 11575 39899
rect 16298 39896 16304 39908
rect 15686 39868 16304 39896
rect 11517 39859 11575 39865
rect 16298 39856 16304 39868
rect 16356 39896 16362 39908
rect 18322 39896 18328 39908
rect 16356 39868 16790 39896
rect 17696 39868 18328 39896
rect 16356 39856 16362 39868
rect 11149 39831 11207 39837
rect 11149 39797 11161 39831
rect 11195 39797 11207 39831
rect 11149 39791 11207 39797
rect 11606 39788 11612 39840
rect 11664 39788 11670 39840
rect 12618 39788 12624 39840
rect 12676 39788 12682 39840
rect 15933 39831 15991 39837
rect 15933 39797 15945 39831
rect 15979 39828 15991 39831
rect 17696 39828 17724 39868
rect 18322 39856 18328 39868
rect 18380 39856 18386 39908
rect 19886 39856 19892 39908
rect 19944 39856 19950 39908
rect 21361 39899 21419 39905
rect 21361 39896 21373 39899
rect 20180 39868 21373 39896
rect 15979 39800 17724 39828
rect 17957 39831 18015 39837
rect 15979 39797 15991 39800
rect 15933 39791 15991 39797
rect 17957 39797 17969 39831
rect 18003 39828 18015 39831
rect 18046 39828 18052 39840
rect 18003 39800 18052 39828
rect 18003 39797 18015 39800
rect 17957 39791 18015 39797
rect 18046 39788 18052 39800
rect 18104 39828 18110 39840
rect 18506 39828 18512 39840
rect 18104 39800 18512 39828
rect 18104 39788 18110 39800
rect 18506 39788 18512 39800
rect 18564 39788 18570 39840
rect 19058 39788 19064 39840
rect 19116 39788 19122 39840
rect 19150 39788 19156 39840
rect 19208 39828 19214 39840
rect 20180 39828 20208 39868
rect 21361 39865 21373 39868
rect 21407 39865 21419 39899
rect 21361 39859 21419 39865
rect 22465 39899 22523 39905
rect 22465 39865 22477 39899
rect 22511 39896 22523 39899
rect 24946 39896 24952 39908
rect 22511 39868 24952 39896
rect 22511 39865 22523 39868
rect 22465 39859 22523 39865
rect 24946 39856 24952 39868
rect 25004 39856 25010 39908
rect 19208 39800 20208 39828
rect 19208 39788 19214 39800
rect 22738 39788 22744 39840
rect 22796 39828 22802 39840
rect 22925 39831 22983 39837
rect 22925 39828 22937 39831
rect 22796 39800 22937 39828
rect 22796 39788 22802 39800
rect 22925 39797 22937 39800
rect 22971 39797 22983 39831
rect 22925 39791 22983 39797
rect 23385 39831 23443 39837
rect 23385 39797 23397 39831
rect 23431 39828 23443 39831
rect 24670 39828 24676 39840
rect 23431 39800 24676 39828
rect 23431 39797 23443 39800
rect 23385 39791 23443 39797
rect 24670 39788 24676 39800
rect 24728 39788 24734 39840
rect 25225 39831 25283 39837
rect 25225 39797 25237 39831
rect 25271 39828 25283 39831
rect 26050 39828 26056 39840
rect 25271 39800 26056 39828
rect 25271 39797 25283 39800
rect 25225 39791 25283 39797
rect 26050 39788 26056 39800
rect 26108 39788 26114 39840
rect 26988 39828 27016 39927
rect 39022 39924 39028 39936
rect 39080 39924 39086 39976
rect 39132 39964 39160 39995
rect 39482 39992 39488 40044
rect 39540 39992 39546 40044
rect 40126 39992 40132 40044
rect 40184 39992 40190 40044
rect 40218 39992 40224 40044
rect 40276 40032 40282 40044
rect 43070 40032 43076 40044
rect 40276 40004 43076 40032
rect 40276 39992 40282 40004
rect 40880 39976 40908 40004
rect 43070 39992 43076 40004
rect 43128 39992 43134 40044
rect 43714 39992 43720 40044
rect 43772 40032 43778 40044
rect 43993 40035 44051 40041
rect 43993 40032 44005 40035
rect 43772 40004 44005 40032
rect 43772 39992 43778 40004
rect 43993 40001 44005 40004
rect 44039 40001 44051 40035
rect 43993 39995 44051 40001
rect 44082 39992 44088 40044
rect 44140 40032 44146 40044
rect 44192 40041 44220 40072
rect 44177 40035 44235 40041
rect 44177 40032 44189 40035
rect 44140 40004 44189 40032
rect 44140 39992 44146 40004
rect 44177 40001 44189 40004
rect 44223 40001 44235 40035
rect 45664 40032 45692 40072
rect 46860 40032 46888 40140
rect 48038 40128 48044 40140
rect 48096 40128 48102 40180
rect 48498 40128 48504 40180
rect 48556 40168 48562 40180
rect 49602 40168 49608 40180
rect 48556 40140 49608 40168
rect 48556 40128 48562 40140
rect 49602 40128 49608 40140
rect 49660 40128 49666 40180
rect 51810 40168 51816 40180
rect 49712 40140 51816 40168
rect 47762 40060 47768 40112
rect 47820 40100 47826 40112
rect 49421 40103 49479 40109
rect 47820 40072 48912 40100
rect 47820 40060 47826 40072
rect 45664 40004 46888 40032
rect 46937 40035 46995 40041
rect 44177 39995 44235 40001
rect 46937 40001 46949 40035
rect 46983 40032 46995 40035
rect 47394 40032 47400 40044
rect 46983 40004 47400 40032
rect 46983 40001 46995 40004
rect 46937 39995 46995 40001
rect 47394 39992 47400 40004
rect 47452 39992 47458 40044
rect 48884 40041 48912 40072
rect 49421 40069 49433 40103
rect 49467 40069 49479 40103
rect 49421 40063 49479 40069
rect 48869 40035 48927 40041
rect 48869 40001 48881 40035
rect 48915 40032 48927 40035
rect 49436 40032 49464 40063
rect 49510 40060 49516 40112
rect 49568 40100 49574 40112
rect 49712 40100 49740 40140
rect 51810 40128 51816 40140
rect 51868 40128 51874 40180
rect 56321 40171 56379 40177
rect 56321 40137 56333 40171
rect 56367 40168 56379 40171
rect 56594 40168 56600 40180
rect 56367 40140 56600 40168
rect 56367 40137 56379 40140
rect 56321 40131 56379 40137
rect 56594 40128 56600 40140
rect 56652 40128 56658 40180
rect 57514 40128 57520 40180
rect 57572 40168 57578 40180
rect 57572 40140 58848 40168
rect 57572 40128 57578 40140
rect 49568 40072 49740 40100
rect 49568 40060 49574 40072
rect 57146 40060 57152 40112
rect 57204 40100 57210 40112
rect 58710 40100 58716 40112
rect 57204 40072 58716 40100
rect 57204 40060 57210 40072
rect 51077 40035 51135 40041
rect 51077 40032 51089 40035
rect 48915 40004 49280 40032
rect 49436 40004 51089 40032
rect 48915 40001 48927 40004
rect 48869 39995 48927 40001
rect 39669 39967 39727 39973
rect 39669 39964 39681 39967
rect 39132 39936 39681 39964
rect 39669 39933 39681 39936
rect 39715 39964 39727 39967
rect 40681 39967 40739 39973
rect 40681 39964 40693 39967
rect 39715 39936 40693 39964
rect 39715 39933 39727 39936
rect 39669 39927 39727 39933
rect 40681 39933 40693 39936
rect 40727 39933 40739 39967
rect 40681 39927 40739 39933
rect 40862 39924 40868 39976
rect 40920 39924 40926 39976
rect 42426 39924 42432 39976
rect 42484 39964 42490 39976
rect 45370 39964 45376 39976
rect 42484 39936 45376 39964
rect 42484 39924 42490 39936
rect 45370 39924 45376 39936
rect 45428 39924 45434 39976
rect 47121 39967 47179 39973
rect 47121 39933 47133 39967
rect 47167 39933 47179 39967
rect 47121 39927 47179 39933
rect 48041 39967 48099 39973
rect 48041 39933 48053 39967
rect 48087 39964 48099 39967
rect 48406 39964 48412 39976
rect 48087 39936 48412 39964
rect 48087 39933 48099 39936
rect 48041 39927 48099 39933
rect 27338 39856 27344 39908
rect 27396 39856 27402 39908
rect 28626 39896 28632 39908
rect 28566 39868 28632 39896
rect 28626 39856 28632 39868
rect 28684 39856 28690 39908
rect 29365 39899 29423 39905
rect 29365 39865 29377 39899
rect 29411 39896 29423 39899
rect 29822 39896 29828 39908
rect 29411 39868 29828 39896
rect 29411 39865 29423 39868
rect 29365 39859 29423 39865
rect 29822 39856 29828 39868
rect 29880 39856 29886 39908
rect 30101 39899 30159 39905
rect 30101 39865 30113 39899
rect 30147 39896 30159 39899
rect 30374 39896 30380 39908
rect 30147 39868 30380 39896
rect 30147 39865 30159 39868
rect 30101 39859 30159 39865
rect 30374 39856 30380 39868
rect 30432 39856 30438 39908
rect 30558 39856 30564 39908
rect 30616 39856 30622 39908
rect 32582 39856 32588 39908
rect 32640 39896 32646 39908
rect 33318 39896 33324 39908
rect 32640 39868 33324 39896
rect 32640 39856 32646 39868
rect 33318 39856 33324 39868
rect 33376 39896 33382 39908
rect 35526 39896 35532 39908
rect 33376 39868 35532 39896
rect 33376 39856 33382 39868
rect 35526 39856 35532 39868
rect 35584 39896 35590 39908
rect 35584 39868 35650 39896
rect 35584 39856 35590 39868
rect 36814 39856 36820 39908
rect 36872 39856 36878 39908
rect 41141 39899 41199 39905
rect 38948 39868 40172 39896
rect 27430 39828 27436 39840
rect 26988 39800 27436 39828
rect 27430 39788 27436 39800
rect 27488 39788 27494 39840
rect 28902 39788 28908 39840
rect 28960 39828 28966 39840
rect 28997 39831 29055 39837
rect 28997 39828 29009 39831
rect 28960 39800 29009 39828
rect 28960 39788 28966 39800
rect 28997 39797 29009 39800
rect 29043 39797 29055 39831
rect 28997 39791 29055 39797
rect 29457 39831 29515 39837
rect 29457 39797 29469 39831
rect 29503 39828 29515 39831
rect 30742 39828 30748 39840
rect 29503 39800 30748 39828
rect 29503 39797 29515 39800
rect 29457 39791 29515 39797
rect 30742 39788 30748 39800
rect 30800 39788 30806 39840
rect 31570 39788 31576 39840
rect 31628 39788 31634 39840
rect 32950 39788 32956 39840
rect 33008 39788 33014 39840
rect 35250 39788 35256 39840
rect 35308 39828 35314 39840
rect 35345 39831 35403 39837
rect 35345 39828 35357 39831
rect 35308 39800 35357 39828
rect 35308 39788 35314 39800
rect 35345 39797 35357 39800
rect 35391 39828 35403 39831
rect 35986 39828 35992 39840
rect 35391 39800 35992 39828
rect 35391 39797 35403 39800
rect 35345 39791 35403 39797
rect 35986 39788 35992 39800
rect 36044 39788 36050 39840
rect 37274 39788 37280 39840
rect 37332 39828 37338 39840
rect 38948 39828 38976 39868
rect 37332 39800 38976 39828
rect 37332 39788 37338 39800
rect 39022 39788 39028 39840
rect 39080 39828 39086 39840
rect 39390 39828 39396 39840
rect 39080 39800 39396 39828
rect 39080 39788 39086 39800
rect 39390 39788 39396 39800
rect 39448 39788 39454 39840
rect 39577 39831 39635 39837
rect 39577 39797 39589 39831
rect 39623 39828 39635 39831
rect 39666 39828 39672 39840
rect 39623 39800 39672 39828
rect 39623 39797 39635 39800
rect 39577 39791 39635 39797
rect 39666 39788 39672 39800
rect 39724 39788 39730 39840
rect 39850 39788 39856 39840
rect 39908 39828 39914 39840
rect 40037 39831 40095 39837
rect 40037 39828 40049 39831
rect 39908 39800 40049 39828
rect 39908 39788 39914 39800
rect 40037 39797 40049 39800
rect 40083 39797 40095 39831
rect 40144 39828 40172 39868
rect 41141 39865 41153 39899
rect 41187 39896 41199 39899
rect 41414 39896 41420 39908
rect 41187 39868 41420 39896
rect 41187 39865 41199 39868
rect 41141 39859 41199 39865
rect 41414 39856 41420 39868
rect 41472 39856 41478 39908
rect 41874 39856 41880 39908
rect 41932 39856 41938 39908
rect 43349 39899 43407 39905
rect 43349 39896 43361 39899
rect 42536 39868 43361 39896
rect 42536 39828 42564 39868
rect 43349 39865 43361 39868
rect 43395 39896 43407 39899
rect 43901 39899 43959 39905
rect 43901 39896 43913 39899
rect 43395 39868 43913 39896
rect 43395 39865 43407 39868
rect 43349 39859 43407 39865
rect 43901 39865 43913 39868
rect 43947 39865 43959 39899
rect 43901 39859 43959 39865
rect 46198 39856 46204 39908
rect 46256 39896 46262 39908
rect 46256 39868 46612 39896
rect 46256 39856 46262 39868
rect 40144 39800 42564 39828
rect 42613 39831 42671 39837
rect 40037 39791 40095 39797
rect 42613 39797 42625 39831
rect 42659 39828 42671 39831
rect 42886 39828 42892 39840
rect 42659 39800 42892 39828
rect 42659 39797 42671 39800
rect 42613 39791 42671 39797
rect 42886 39788 42892 39800
rect 42944 39828 42950 39840
rect 43254 39828 43260 39840
rect 42944 39800 43260 39828
rect 42944 39788 42950 39800
rect 43254 39788 43260 39800
rect 43312 39788 43318 39840
rect 43530 39788 43536 39840
rect 43588 39788 43594 39840
rect 45186 39788 45192 39840
rect 45244 39828 45250 39840
rect 46474 39828 46480 39840
rect 45244 39800 46480 39828
rect 45244 39788 45250 39800
rect 46474 39788 46480 39800
rect 46532 39788 46538 39840
rect 46584 39828 46612 39868
rect 46658 39856 46664 39908
rect 46716 39896 46722 39908
rect 47136 39896 47164 39927
rect 48406 39924 48412 39936
rect 48464 39924 48470 39976
rect 49050 39924 49056 39976
rect 49108 39924 49114 39976
rect 49252 39896 49280 40004
rect 51077 40001 51089 40004
rect 51123 40001 51135 40035
rect 51077 39995 51135 40001
rect 51353 40035 51411 40041
rect 51353 40001 51365 40035
rect 51399 40032 51411 40035
rect 52454 40032 52460 40044
rect 51399 40004 52460 40032
rect 51399 40001 51411 40004
rect 51353 39995 51411 40001
rect 52454 39992 52460 40004
rect 52512 39992 52518 40044
rect 53650 39992 53656 40044
rect 53708 40032 53714 40044
rect 55674 40032 55680 40044
rect 53708 40004 55680 40032
rect 53708 39992 53714 40004
rect 55674 39992 55680 40004
rect 55732 39992 55738 40044
rect 57808 40041 57836 40072
rect 58710 40060 58716 40072
rect 58768 40060 58774 40112
rect 57793 40035 57851 40041
rect 57793 40001 57805 40035
rect 57839 40001 57851 40035
rect 57793 39995 57851 40001
rect 58621 40035 58679 40041
rect 58621 40001 58633 40035
rect 58667 40032 58679 40035
rect 58820 40032 58848 40140
rect 58667 40004 58848 40032
rect 58667 40001 58679 40004
rect 58621 39995 58679 40001
rect 49970 39924 49976 39976
rect 50028 39924 50034 39976
rect 51997 39967 52055 39973
rect 51997 39933 52009 39967
rect 52043 39964 52055 39967
rect 53742 39964 53748 39976
rect 52043 39936 53748 39964
rect 52043 39933 52055 39936
rect 51997 39927 52055 39933
rect 49786 39896 49792 39908
rect 46716 39868 47164 39896
rect 47228 39868 49096 39896
rect 49252 39868 49792 39896
rect 46716 39856 46722 39868
rect 47228 39828 47256 39868
rect 46584 39800 47256 39828
rect 47394 39788 47400 39840
rect 47452 39828 47458 39840
rect 47765 39831 47823 39837
rect 47765 39828 47777 39831
rect 47452 39800 47777 39828
rect 47452 39788 47458 39800
rect 47765 39797 47777 39800
rect 47811 39797 47823 39831
rect 47765 39791 47823 39797
rect 48590 39788 48596 39840
rect 48648 39788 48654 39840
rect 48958 39788 48964 39840
rect 49016 39788 49022 39840
rect 49068 39828 49096 39868
rect 49786 39856 49792 39868
rect 49844 39856 49850 39908
rect 49988 39828 50016 39924
rect 49068 39800 50016 39828
rect 50154 39788 50160 39840
rect 50212 39828 50218 39840
rect 50890 39828 50896 39840
rect 50212 39800 50896 39828
rect 50212 39788 50218 39800
rect 50890 39788 50896 39800
rect 50948 39828 50954 39840
rect 52012 39828 52040 39927
rect 53742 39924 53748 39936
rect 53800 39924 53806 39976
rect 57698 39924 57704 39976
rect 57756 39924 57762 39976
rect 52822 39856 52828 39908
rect 52880 39896 52886 39908
rect 55306 39896 55312 39908
rect 52880 39868 55312 39896
rect 52880 39856 52886 39868
rect 55306 39856 55312 39868
rect 55364 39896 55370 39908
rect 55861 39899 55919 39905
rect 55861 39896 55873 39899
rect 55364 39868 55873 39896
rect 55364 39856 55370 39868
rect 55861 39865 55873 39868
rect 55907 39865 55919 39899
rect 55861 39859 55919 39865
rect 56965 39899 57023 39905
rect 56965 39865 56977 39899
rect 57011 39896 57023 39899
rect 57330 39896 57336 39908
rect 57011 39868 57336 39896
rect 57011 39865 57023 39868
rect 56965 39859 57023 39865
rect 57330 39856 57336 39868
rect 57388 39856 57394 39908
rect 57609 39899 57667 39905
rect 57609 39865 57621 39899
rect 57655 39896 57667 39899
rect 58802 39896 58808 39908
rect 57655 39868 58808 39896
rect 57655 39865 57667 39868
rect 57609 39859 57667 39865
rect 58802 39856 58808 39868
rect 58860 39856 58866 39908
rect 50948 39800 52040 39828
rect 50948 39788 50954 39800
rect 55214 39788 55220 39840
rect 55272 39828 55278 39840
rect 55401 39831 55459 39837
rect 55401 39828 55413 39831
rect 55272 39800 55413 39828
rect 55272 39788 55278 39800
rect 55401 39797 55413 39800
rect 55447 39828 55459 39831
rect 55766 39828 55772 39840
rect 55447 39800 55772 39828
rect 55447 39797 55459 39800
rect 55401 39791 55459 39797
rect 55766 39788 55772 39800
rect 55824 39828 55830 39840
rect 55953 39831 56011 39837
rect 55953 39828 55965 39831
rect 55824 39800 55965 39828
rect 55824 39788 55830 39800
rect 55953 39797 55965 39800
rect 55999 39797 56011 39831
rect 55953 39791 56011 39797
rect 57238 39788 57244 39840
rect 57296 39788 57302 39840
rect 58066 39788 58072 39840
rect 58124 39788 58130 39840
rect 58434 39788 58440 39840
rect 58492 39788 58498 39840
rect 58529 39831 58587 39837
rect 58529 39797 58541 39831
rect 58575 39828 58587 39831
rect 58894 39828 58900 39840
rect 58575 39800 58900 39828
rect 58575 39797 58587 39800
rect 58529 39791 58587 39797
rect 58894 39788 58900 39800
rect 58952 39788 58958 39840
rect 552 39738 66424 39760
rect 552 39686 2918 39738
rect 2970 39686 2982 39738
rect 3034 39686 3046 39738
rect 3098 39686 3110 39738
rect 3162 39686 3174 39738
rect 3226 39686 51918 39738
rect 51970 39686 51982 39738
rect 52034 39686 52046 39738
rect 52098 39686 52110 39738
rect 52162 39686 52174 39738
rect 52226 39686 66424 39738
rect 552 39664 66424 39686
rect 14182 39624 14188 39636
rect 10428 39596 14188 39624
rect 9674 39516 9680 39568
rect 9732 39516 9738 39568
rect 10134 39516 10140 39568
rect 10192 39516 10198 39568
rect 10428 39497 10456 39596
rect 14182 39584 14188 39596
rect 14240 39584 14246 39636
rect 15197 39627 15255 39633
rect 15197 39593 15209 39627
rect 15243 39624 15255 39627
rect 15286 39624 15292 39636
rect 15243 39596 15292 39624
rect 15243 39593 15255 39596
rect 15197 39587 15255 39593
rect 15286 39584 15292 39596
rect 15344 39584 15350 39636
rect 15562 39584 15568 39636
rect 15620 39584 15626 39636
rect 15657 39627 15715 39633
rect 15657 39593 15669 39627
rect 15703 39624 15715 39627
rect 16301 39627 16359 39633
rect 16301 39624 16313 39627
rect 15703 39596 16313 39624
rect 15703 39593 15715 39596
rect 15657 39587 15715 39593
rect 16301 39593 16313 39596
rect 16347 39593 16359 39627
rect 16301 39587 16359 39593
rect 16482 39584 16488 39636
rect 16540 39624 16546 39636
rect 16761 39627 16819 39633
rect 16761 39624 16773 39627
rect 16540 39596 16773 39624
rect 16540 39584 16546 39596
rect 16761 39593 16773 39596
rect 16807 39593 16819 39627
rect 16761 39587 16819 39593
rect 17954 39584 17960 39636
rect 18012 39624 18018 39636
rect 18233 39627 18291 39633
rect 18233 39624 18245 39627
rect 18012 39596 18245 39624
rect 18012 39584 18018 39596
rect 18233 39593 18245 39596
rect 18279 39593 18291 39627
rect 18233 39587 18291 39593
rect 18693 39627 18751 39633
rect 18693 39593 18705 39627
rect 18739 39624 18751 39627
rect 19150 39624 19156 39636
rect 18739 39596 19156 39624
rect 18739 39593 18751 39596
rect 18693 39587 18751 39593
rect 19150 39584 19156 39596
rect 19208 39584 19214 39636
rect 20070 39584 20076 39636
rect 20128 39624 20134 39636
rect 21542 39624 21548 39636
rect 20128 39596 21548 39624
rect 20128 39584 20134 39596
rect 21542 39584 21548 39596
rect 21600 39624 21606 39636
rect 21600 39596 24532 39624
rect 21600 39584 21606 39596
rect 12894 39516 12900 39568
rect 12952 39516 12958 39568
rect 14461 39559 14519 39565
rect 14461 39525 14473 39559
rect 14507 39556 14519 39559
rect 14550 39556 14556 39568
rect 14507 39528 14556 39556
rect 14507 39525 14519 39528
rect 14461 39519 14519 39525
rect 14550 39516 14556 39528
rect 14608 39516 14614 39568
rect 16209 39559 16267 39565
rect 16209 39525 16221 39559
rect 16255 39556 16267 39559
rect 16669 39559 16727 39565
rect 16669 39556 16681 39559
rect 16255 39528 16681 39556
rect 16255 39525 16267 39528
rect 16209 39519 16267 39525
rect 16669 39525 16681 39528
rect 16715 39556 16727 39559
rect 17770 39556 17776 39568
rect 16715 39528 17776 39556
rect 16715 39525 16727 39528
rect 16669 39519 16727 39525
rect 17770 39516 17776 39528
rect 17828 39516 17834 39568
rect 18782 39516 18788 39568
rect 18840 39516 18846 39568
rect 19058 39516 19064 39568
rect 19116 39556 19122 39568
rect 21729 39559 21787 39565
rect 21729 39556 21741 39559
rect 19116 39528 21741 39556
rect 19116 39516 19122 39528
rect 21729 39525 21741 39528
rect 21775 39525 21787 39559
rect 21729 39519 21787 39525
rect 10413 39491 10471 39497
rect 10413 39457 10425 39491
rect 10459 39457 10471 39491
rect 10413 39451 10471 39457
rect 11330 39448 11336 39500
rect 11388 39448 11394 39500
rect 11425 39491 11483 39497
rect 11425 39457 11437 39491
rect 11471 39488 11483 39491
rect 12066 39488 12072 39500
rect 11471 39460 12072 39488
rect 11471 39457 11483 39460
rect 11425 39451 11483 39457
rect 12066 39448 12072 39460
rect 12124 39448 12130 39500
rect 14369 39491 14427 39497
rect 14369 39457 14381 39491
rect 14415 39488 14427 39491
rect 15102 39488 15108 39500
rect 14415 39460 15108 39488
rect 14415 39457 14427 39460
rect 14369 39451 14427 39457
rect 15102 39448 15108 39460
rect 15160 39448 15166 39500
rect 17494 39448 17500 39500
rect 17552 39448 17558 39500
rect 17589 39491 17647 39497
rect 17589 39457 17601 39491
rect 17635 39488 17647 39491
rect 18046 39488 18052 39500
rect 17635 39460 18052 39488
rect 17635 39457 17647 39460
rect 17589 39451 17647 39457
rect 18046 39448 18052 39460
rect 18104 39448 18110 39500
rect 18325 39491 18383 39497
rect 18325 39457 18337 39491
rect 18371 39488 18383 39491
rect 20622 39488 20628 39500
rect 18371 39460 20628 39488
rect 18371 39457 18383 39460
rect 18325 39451 18383 39457
rect 20622 39448 20628 39460
rect 20680 39448 20686 39500
rect 21634 39448 21640 39500
rect 21692 39448 21698 39500
rect 22480 39497 22508 39596
rect 22738 39516 22744 39568
rect 22796 39516 22802 39568
rect 24504 39497 24532 39596
rect 25038 39584 25044 39636
rect 25096 39624 25102 39636
rect 25590 39624 25596 39636
rect 25096 39596 25596 39624
rect 25096 39584 25102 39596
rect 25590 39584 25596 39596
rect 25648 39624 25654 39636
rect 26142 39624 26148 39636
rect 25648 39596 26148 39624
rect 25648 39584 25654 39596
rect 26142 39584 26148 39596
rect 26200 39584 26206 39636
rect 26234 39584 26240 39636
rect 26292 39584 26298 39636
rect 26418 39584 26424 39636
rect 26476 39584 26482 39636
rect 26510 39584 26516 39636
rect 26568 39624 26574 39636
rect 26881 39627 26939 39633
rect 26881 39624 26893 39627
rect 26568 39596 26893 39624
rect 26568 39584 26574 39596
rect 26881 39593 26893 39596
rect 26927 39624 26939 39627
rect 26970 39624 26976 39636
rect 26927 39596 26976 39624
rect 26927 39593 26939 39596
rect 26881 39587 26939 39593
rect 26970 39584 26976 39596
rect 27028 39584 27034 39636
rect 27338 39584 27344 39636
rect 27396 39624 27402 39636
rect 27709 39627 27767 39633
rect 27709 39624 27721 39627
rect 27396 39596 27721 39624
rect 27396 39584 27402 39596
rect 27709 39593 27721 39596
rect 27755 39593 27767 39627
rect 27709 39587 27767 39593
rect 28074 39584 28080 39636
rect 28132 39584 28138 39636
rect 29730 39624 29736 39636
rect 28368 39596 29736 39624
rect 24762 39516 24768 39568
rect 24820 39516 24826 39568
rect 26050 39516 26056 39568
rect 26108 39556 26114 39568
rect 26789 39559 26847 39565
rect 26789 39556 26801 39559
rect 26108 39528 26801 39556
rect 26108 39516 26114 39528
rect 26789 39525 26801 39528
rect 26835 39556 26847 39559
rect 27614 39556 27620 39568
rect 26835 39528 27620 39556
rect 26835 39525 26847 39528
rect 26789 39519 26847 39525
rect 27614 39516 27620 39528
rect 27672 39516 27678 39568
rect 22465 39491 22523 39497
rect 22465 39457 22477 39491
rect 22511 39457 22523 39491
rect 24489 39491 24547 39497
rect 23874 39460 24440 39488
rect 22465 39451 22523 39457
rect 8202 39380 8208 39432
rect 8260 39420 8266 39432
rect 8389 39423 8447 39429
rect 8389 39420 8401 39423
rect 8260 39392 8401 39420
rect 8260 39380 8266 39392
rect 8389 39389 8401 39392
rect 8435 39389 8447 39423
rect 8389 39383 8447 39389
rect 8665 39423 8723 39429
rect 8665 39389 8677 39423
rect 8711 39420 8723 39423
rect 11348 39420 11376 39448
rect 8711 39392 11376 39420
rect 8711 39389 8723 39392
rect 8665 39383 8723 39389
rect 11606 39380 11612 39432
rect 11664 39380 11670 39432
rect 12161 39423 12219 39429
rect 12161 39389 12173 39423
rect 12207 39389 12219 39423
rect 12161 39383 12219 39389
rect 12437 39423 12495 39429
rect 12437 39389 12449 39423
rect 12483 39420 12495 39423
rect 12526 39420 12532 39432
rect 12483 39392 12532 39420
rect 12483 39389 12495 39392
rect 12437 39383 12495 39389
rect 10410 39312 10416 39364
rect 10468 39352 10474 39364
rect 11624 39352 11652 39380
rect 10468 39324 11652 39352
rect 10468 39312 10474 39324
rect 7834 39244 7840 39296
rect 7892 39244 7898 39296
rect 10318 39244 10324 39296
rect 10376 39284 10382 39296
rect 10965 39287 11023 39293
rect 10965 39284 10977 39287
rect 10376 39256 10977 39284
rect 10376 39244 10382 39256
rect 10965 39253 10977 39256
rect 11011 39253 11023 39287
rect 12176 39284 12204 39383
rect 12526 39380 12532 39392
rect 12584 39380 12590 39432
rect 14553 39423 14611 39429
rect 14553 39389 14565 39423
rect 14599 39389 14611 39423
rect 14553 39383 14611 39389
rect 15841 39423 15899 39429
rect 15841 39389 15853 39423
rect 15887 39420 15899 39423
rect 16758 39420 16764 39432
rect 15887 39392 16764 39420
rect 15887 39389 15899 39392
rect 15841 39383 15899 39389
rect 13814 39312 13820 39364
rect 13872 39352 13878 39364
rect 14568 39352 14596 39383
rect 16758 39380 16764 39392
rect 16816 39380 16822 39432
rect 16945 39423 17003 39429
rect 16945 39389 16957 39423
rect 16991 39420 17003 39423
rect 17310 39420 17316 39432
rect 16991 39392 17316 39420
rect 16991 39389 17003 39392
rect 16945 39383 17003 39389
rect 17310 39380 17316 39392
rect 17368 39380 17374 39432
rect 17773 39423 17831 39429
rect 17773 39389 17785 39423
rect 17819 39389 17831 39423
rect 17773 39383 17831 39389
rect 18141 39423 18199 39429
rect 18141 39389 18153 39423
rect 18187 39389 18199 39423
rect 18141 39383 18199 39389
rect 15378 39352 15384 39364
rect 13872 39324 15384 39352
rect 13872 39312 13878 39324
rect 15378 39312 15384 39324
rect 15436 39312 15442 39364
rect 12434 39284 12440 39296
rect 12176 39256 12440 39284
rect 10965 39247 11023 39253
rect 12434 39244 12440 39256
rect 12492 39284 12498 39296
rect 13538 39284 13544 39296
rect 12492 39256 13544 39284
rect 12492 39244 12498 39256
rect 13538 39244 13544 39256
rect 13596 39244 13602 39296
rect 13906 39244 13912 39296
rect 13964 39244 13970 39296
rect 13998 39244 14004 39296
rect 14056 39244 14062 39296
rect 16850 39244 16856 39296
rect 16908 39284 16914 39296
rect 17129 39287 17187 39293
rect 17129 39284 17141 39287
rect 16908 39256 17141 39284
rect 16908 39244 16914 39256
rect 17129 39253 17141 39256
rect 17175 39253 17187 39287
rect 17788 39284 17816 39383
rect 18156 39352 18184 39383
rect 18874 39380 18880 39432
rect 18932 39420 18938 39432
rect 21358 39420 21364 39432
rect 18932 39392 21364 39420
rect 18932 39380 18938 39392
rect 21358 39380 21364 39392
rect 21416 39380 21422 39432
rect 21818 39380 21824 39432
rect 21876 39380 21882 39432
rect 24210 39380 24216 39432
rect 24268 39380 24274 39432
rect 24412 39420 24440 39460
rect 24489 39457 24501 39491
rect 24535 39457 24547 39491
rect 24489 39451 24547 39457
rect 25222 39420 25228 39432
rect 24412 39392 25228 39420
rect 25222 39380 25228 39392
rect 25280 39420 25286 39432
rect 25884 39420 25912 39474
rect 26234 39448 26240 39500
rect 26292 39488 26298 39500
rect 27246 39488 27252 39500
rect 26292 39460 27252 39488
rect 26292 39448 26298 39460
rect 25280 39392 25912 39420
rect 25280 39380 25286 39392
rect 26142 39380 26148 39432
rect 26200 39420 26206 39432
rect 26510 39420 26516 39432
rect 26200 39392 26516 39420
rect 26200 39380 26206 39392
rect 26510 39380 26516 39392
rect 26568 39380 26574 39432
rect 26988 39429 27016 39460
rect 27246 39448 27252 39460
rect 27304 39448 27310 39500
rect 27430 39448 27436 39500
rect 27488 39448 27494 39500
rect 26973 39423 27031 39429
rect 26973 39389 26985 39423
rect 27019 39389 27031 39423
rect 26973 39383 27031 39389
rect 28166 39380 28172 39432
rect 28224 39380 28230 39432
rect 28261 39423 28319 39429
rect 28261 39389 28273 39423
rect 28307 39389 28319 39423
rect 28261 39383 28319 39389
rect 18414 39352 18420 39364
rect 18156 39324 18420 39352
rect 18414 39312 18420 39324
rect 18472 39312 18478 39364
rect 19978 39352 19984 39364
rect 19812 39324 19984 39352
rect 19812 39284 19840 39324
rect 19978 39312 19984 39324
rect 20036 39352 20042 39364
rect 20622 39352 20628 39364
rect 20036 39324 20628 39352
rect 20036 39312 20042 39324
rect 20622 39312 20628 39324
rect 20680 39312 20686 39364
rect 20806 39312 20812 39364
rect 20864 39352 20870 39364
rect 20864 39324 22094 39352
rect 20864 39312 20870 39324
rect 17788 39256 19840 39284
rect 17129 39247 17187 39253
rect 19886 39244 19892 39296
rect 19944 39284 19950 39296
rect 21269 39287 21327 39293
rect 21269 39284 21281 39287
rect 19944 39256 21281 39284
rect 19944 39244 19950 39256
rect 21269 39253 21281 39256
rect 21315 39253 21327 39287
rect 22066 39284 22094 39324
rect 26786 39312 26792 39364
rect 26844 39352 26850 39364
rect 28276 39352 28304 39383
rect 26844 39324 28304 39352
rect 26844 39312 26850 39324
rect 28368 39284 28396 39596
rect 29730 39584 29736 39596
rect 29788 39584 29794 39636
rect 30374 39584 30380 39636
rect 30432 39584 30438 39636
rect 31294 39584 31300 39636
rect 31352 39624 31358 39636
rect 32582 39624 32588 39636
rect 31352 39596 32588 39624
rect 31352 39584 31358 39596
rect 32582 39584 32588 39596
rect 32640 39584 32646 39636
rect 33134 39584 33140 39636
rect 33192 39624 33198 39636
rect 33781 39627 33839 39633
rect 33781 39624 33793 39627
rect 33192 39596 33793 39624
rect 33192 39584 33198 39596
rect 33781 39593 33793 39596
rect 33827 39593 33839 39627
rect 33781 39587 33839 39593
rect 33962 39584 33968 39636
rect 34020 39624 34026 39636
rect 34020 39596 34560 39624
rect 34020 39584 34026 39596
rect 28813 39559 28871 39565
rect 28813 39525 28825 39559
rect 28859 39556 28871 39559
rect 28902 39556 28908 39568
rect 28859 39528 28908 39556
rect 28859 39525 28871 39528
rect 28813 39519 28871 39525
rect 28902 39516 28908 39528
rect 28960 39516 28966 39568
rect 30098 39516 30104 39568
rect 30156 39556 30162 39568
rect 30156 39528 31984 39556
rect 30156 39516 30162 39528
rect 31956 39500 31984 39528
rect 32122 39516 32128 39568
rect 32180 39556 32186 39568
rect 32217 39559 32275 39565
rect 32217 39556 32229 39559
rect 32180 39528 32229 39556
rect 32180 39516 32186 39528
rect 32217 39525 32229 39528
rect 32263 39525 32275 39559
rect 32600 39556 32628 39584
rect 32600 39528 32706 39556
rect 32217 39519 32275 39525
rect 29914 39448 29920 39500
rect 29972 39448 29978 39500
rect 30208 39460 30420 39488
rect 28537 39423 28595 39429
rect 28537 39389 28549 39423
rect 28583 39420 28595 39423
rect 28583 39392 28672 39420
rect 28583 39389 28595 39392
rect 28537 39383 28595 39389
rect 22066 39256 28396 39284
rect 28644 39284 28672 39392
rect 28810 39380 28816 39432
rect 28868 39420 28874 39432
rect 30208 39420 30236 39460
rect 28868 39392 30236 39420
rect 30392 39420 30420 39460
rect 30466 39448 30472 39500
rect 30524 39488 30530 39500
rect 30745 39491 30803 39497
rect 30745 39488 30757 39491
rect 30524 39460 30757 39488
rect 30524 39448 30530 39460
rect 30745 39457 30757 39460
rect 30791 39457 30803 39491
rect 30745 39451 30803 39457
rect 31938 39448 31944 39500
rect 31996 39448 32002 39500
rect 34330 39448 34336 39500
rect 34388 39448 34394 39500
rect 34532 39488 34560 39596
rect 35434 39584 35440 39636
rect 35492 39624 35498 39636
rect 35621 39627 35679 39633
rect 35621 39624 35633 39627
rect 35492 39596 35633 39624
rect 35492 39584 35498 39596
rect 35621 39593 35633 39596
rect 35667 39593 35679 39627
rect 35621 39587 35679 39593
rect 36725 39627 36783 39633
rect 36725 39593 36737 39627
rect 36771 39624 36783 39627
rect 36814 39624 36820 39636
rect 36771 39596 36820 39624
rect 36771 39593 36783 39596
rect 36725 39587 36783 39593
rect 36814 39584 36820 39596
rect 36872 39584 36878 39636
rect 36906 39584 36912 39636
rect 36964 39624 36970 39636
rect 38381 39627 38439 39633
rect 38381 39624 38393 39627
rect 36964 39596 38393 39624
rect 36964 39584 36970 39596
rect 38381 39593 38393 39596
rect 38427 39624 38439 39627
rect 39666 39624 39672 39636
rect 38427 39596 39672 39624
rect 38427 39593 38439 39596
rect 38381 39587 38439 39593
rect 39666 39584 39672 39596
rect 39724 39584 39730 39636
rect 40034 39584 40040 39636
rect 40092 39624 40098 39636
rect 40681 39627 40739 39633
rect 40681 39624 40693 39627
rect 40092 39596 40693 39624
rect 40092 39584 40098 39596
rect 40681 39593 40693 39596
rect 40727 39593 40739 39627
rect 40681 39587 40739 39593
rect 40770 39584 40776 39636
rect 40828 39624 40834 39636
rect 40954 39624 40960 39636
rect 40828 39596 40960 39624
rect 40828 39584 40834 39596
rect 40954 39584 40960 39596
rect 41012 39624 41018 39636
rect 42153 39627 42211 39633
rect 42153 39624 42165 39627
rect 41012 39596 42165 39624
rect 41012 39584 41018 39596
rect 42153 39593 42165 39596
rect 42199 39593 42211 39627
rect 42153 39587 42211 39593
rect 42242 39584 42248 39636
rect 42300 39584 42306 39636
rect 43070 39584 43076 39636
rect 43128 39624 43134 39636
rect 43128 39596 44956 39624
rect 43128 39584 43134 39596
rect 35066 39516 35072 39568
rect 35124 39556 35130 39568
rect 36081 39559 36139 39565
rect 36081 39556 36093 39559
rect 35124 39528 36093 39556
rect 35124 39516 35130 39528
rect 36081 39525 36093 39528
rect 36127 39525 36139 39559
rect 36081 39519 36139 39525
rect 36538 39516 36544 39568
rect 36596 39556 36602 39568
rect 37093 39559 37151 39565
rect 37093 39556 37105 39559
rect 36596 39528 37105 39556
rect 36596 39516 36602 39528
rect 37093 39525 37105 39528
rect 37139 39525 37151 39559
rect 37093 39519 37151 39525
rect 39390 39516 39396 39568
rect 39448 39516 39454 39568
rect 39850 39516 39856 39568
rect 39908 39516 39914 39568
rect 43438 39516 43444 39568
rect 43496 39556 43502 39568
rect 43806 39556 43812 39568
rect 43496 39528 43812 39556
rect 43496 39516 43502 39528
rect 43806 39516 43812 39528
rect 43864 39516 43870 39568
rect 34532 39460 35940 39488
rect 30392 39392 30788 39420
rect 28868 39380 28874 39392
rect 30285 39355 30343 39361
rect 30285 39321 30297 39355
rect 30331 39352 30343 39355
rect 30374 39352 30380 39364
rect 30331 39324 30380 39352
rect 30331 39321 30343 39324
rect 30285 39315 30343 39321
rect 30374 39312 30380 39324
rect 30432 39312 30438 39364
rect 30760 39352 30788 39392
rect 30834 39380 30840 39432
rect 30892 39380 30898 39432
rect 31021 39423 31079 39429
rect 31021 39389 31033 39423
rect 31067 39420 31079 39423
rect 31202 39420 31208 39432
rect 31067 39392 31208 39420
rect 31067 39389 31079 39392
rect 31021 39383 31079 39389
rect 31202 39380 31208 39392
rect 31260 39380 31266 39432
rect 34606 39380 34612 39432
rect 34664 39420 34670 39432
rect 34885 39423 34943 39429
rect 34885 39420 34897 39423
rect 34664 39392 34897 39420
rect 34664 39380 34670 39392
rect 34885 39389 34897 39392
rect 34931 39420 34943 39423
rect 35802 39420 35808 39432
rect 34931 39392 35808 39420
rect 34931 39389 34943 39392
rect 34885 39383 34943 39389
rect 35802 39380 35808 39392
rect 35860 39380 35866 39432
rect 35912 39420 35940 39460
rect 35986 39448 35992 39500
rect 36044 39488 36050 39500
rect 38286 39488 38292 39500
rect 36044 39460 36952 39488
rect 36044 39448 36050 39460
rect 36924 39432 36952 39460
rect 37292 39460 38292 39488
rect 36173 39423 36231 39429
rect 36173 39420 36185 39423
rect 35912 39392 36185 39420
rect 36173 39389 36185 39392
rect 36219 39389 36231 39423
rect 36173 39383 36231 39389
rect 36906 39380 36912 39432
rect 36964 39420 36970 39432
rect 37292 39429 37320 39460
rect 38286 39448 38292 39460
rect 38344 39448 38350 39500
rect 40129 39491 40187 39497
rect 40129 39457 40141 39491
rect 40175 39488 40187 39491
rect 40402 39488 40408 39500
rect 40175 39460 40408 39488
rect 40175 39457 40187 39460
rect 40129 39451 40187 39457
rect 40402 39448 40408 39460
rect 40460 39448 40466 39500
rect 40589 39491 40647 39497
rect 40589 39457 40601 39491
rect 40635 39488 40647 39491
rect 41138 39488 41144 39500
rect 40635 39460 41144 39488
rect 40635 39457 40647 39460
rect 40589 39451 40647 39457
rect 41138 39448 41144 39460
rect 41196 39448 41202 39500
rect 41386 39460 42012 39488
rect 37185 39423 37243 39429
rect 37185 39420 37197 39423
rect 36964 39392 37197 39420
rect 36964 39380 36970 39392
rect 37185 39389 37197 39392
rect 37231 39389 37243 39423
rect 37185 39383 37243 39389
rect 37277 39423 37335 39429
rect 37277 39389 37289 39423
rect 37323 39389 37335 39423
rect 37277 39383 37335 39389
rect 37366 39380 37372 39432
rect 37424 39420 37430 39432
rect 37424 39392 40080 39420
rect 37424 39380 37430 39392
rect 40052 39352 40080 39392
rect 40218 39380 40224 39432
rect 40276 39420 40282 39432
rect 40678 39420 40684 39432
rect 40276 39392 40684 39420
rect 40276 39380 40282 39392
rect 40678 39380 40684 39392
rect 40736 39420 40742 39432
rect 40773 39423 40831 39429
rect 40773 39420 40785 39423
rect 40736 39392 40785 39420
rect 40736 39380 40742 39392
rect 40773 39389 40785 39392
rect 40819 39420 40831 39423
rect 41386 39420 41414 39460
rect 40819 39392 41414 39420
rect 40819 39389 40831 39392
rect 40773 39383 40831 39389
rect 41598 39380 41604 39432
rect 41656 39380 41662 39432
rect 41984 39429 42012 39460
rect 43070 39448 43076 39500
rect 43128 39448 43134 39500
rect 44928 39497 44956 39596
rect 45370 39584 45376 39636
rect 45428 39624 45434 39636
rect 45428 39596 46612 39624
rect 45428 39584 45434 39596
rect 46198 39516 46204 39568
rect 46256 39516 46262 39568
rect 44913 39491 44971 39497
rect 44913 39457 44925 39491
rect 44959 39457 44971 39491
rect 46584 39488 46612 39596
rect 46658 39584 46664 39636
rect 46716 39584 46722 39636
rect 47394 39584 47400 39636
rect 47452 39584 47458 39636
rect 48406 39584 48412 39636
rect 48464 39584 48470 39636
rect 48590 39584 48596 39636
rect 48648 39624 48654 39636
rect 48648 39596 49832 39624
rect 48648 39584 48654 39596
rect 49602 39556 49608 39568
rect 49450 39528 49608 39556
rect 49602 39516 49608 39528
rect 49660 39516 49666 39568
rect 49804 39556 49832 39596
rect 50522 39584 50528 39636
rect 50580 39584 50586 39636
rect 50985 39627 51043 39633
rect 50985 39593 50997 39627
rect 51031 39624 51043 39627
rect 51537 39627 51595 39633
rect 51537 39624 51549 39627
rect 51031 39596 51549 39624
rect 51031 39593 51043 39596
rect 50985 39587 51043 39593
rect 51537 39593 51549 39596
rect 51583 39593 51595 39627
rect 51537 39587 51595 39593
rect 54570 39584 54576 39636
rect 54628 39624 54634 39636
rect 54849 39627 54907 39633
rect 54849 39624 54861 39627
rect 54628 39596 54861 39624
rect 54628 39584 54634 39596
rect 54849 39593 54861 39596
rect 54895 39593 54907 39627
rect 54849 39587 54907 39593
rect 54938 39584 54944 39636
rect 54996 39624 55002 39636
rect 55217 39627 55275 39633
rect 55217 39624 55229 39627
rect 54996 39596 55229 39624
rect 54996 39584 55002 39596
rect 55217 39593 55229 39596
rect 55263 39593 55275 39627
rect 55217 39587 55275 39593
rect 55306 39584 55312 39636
rect 55364 39584 55370 39636
rect 55950 39584 55956 39636
rect 56008 39624 56014 39636
rect 56008 39596 57744 39624
rect 56008 39584 56014 39596
rect 51445 39559 51503 39565
rect 51445 39556 51457 39559
rect 49804 39528 51457 39556
rect 51445 39525 51457 39528
rect 51491 39525 51503 39559
rect 51445 39519 51503 39525
rect 53742 39516 53748 39568
rect 53800 39556 53806 39568
rect 56502 39556 56508 39568
rect 53800 39528 56508 39556
rect 53800 39516 53806 39528
rect 56502 39516 56508 39528
rect 56560 39516 56566 39568
rect 57238 39516 57244 39568
rect 57296 39556 57302 39568
rect 57609 39559 57667 39565
rect 57609 39556 57621 39559
rect 57296 39528 57621 39556
rect 57296 39516 57302 39528
rect 57609 39525 57621 39528
rect 57655 39525 57667 39559
rect 57716 39556 57744 39596
rect 58434 39584 58440 39636
rect 58492 39624 58498 39636
rect 59449 39627 59507 39633
rect 59449 39624 59461 39627
rect 58492 39596 59461 39624
rect 58492 39584 58498 39596
rect 59449 39593 59461 39596
rect 59495 39593 59507 39627
rect 59449 39587 59507 39593
rect 57716 39528 58098 39556
rect 57609 39519 57667 39525
rect 46584 39460 48728 39488
rect 44913 39451 44971 39457
rect 41969 39423 42027 39429
rect 41969 39389 41981 39423
rect 42015 39389 42027 39423
rect 41969 39383 42027 39389
rect 43349 39423 43407 39429
rect 43349 39389 43361 39423
rect 43395 39420 43407 39423
rect 43438 39420 43444 39432
rect 43395 39392 43444 39420
rect 43395 39389 43407 39392
rect 43349 39383 43407 39389
rect 43438 39380 43444 39392
rect 43496 39380 43502 39432
rect 43806 39380 43812 39432
rect 43864 39420 43870 39432
rect 44542 39420 44548 39432
rect 43864 39392 44548 39420
rect 43864 39380 43870 39392
rect 44542 39380 44548 39392
rect 44600 39380 44606 39432
rect 45189 39423 45247 39429
rect 45189 39389 45201 39423
rect 45235 39420 45247 39423
rect 45235 39392 47072 39420
rect 45235 39389 45247 39392
rect 45189 39383 45247 39389
rect 47044 39361 47072 39392
rect 47486 39380 47492 39432
rect 47544 39380 47550 39432
rect 47673 39423 47731 39429
rect 47673 39389 47685 39423
rect 47719 39420 47731 39423
rect 47762 39420 47768 39432
rect 47719 39392 47768 39420
rect 47719 39389 47731 39392
rect 47673 39383 47731 39389
rect 47762 39380 47768 39392
rect 47820 39380 47826 39432
rect 48700 39420 48728 39460
rect 50614 39448 50620 39500
rect 50672 39448 50678 39500
rect 50798 39448 50804 39500
rect 50856 39488 50862 39500
rect 52181 39491 52239 39497
rect 50856 39460 51672 39488
rect 50856 39448 50862 39460
rect 49510 39420 49516 39432
rect 48700 39392 49516 39420
rect 49510 39380 49516 39392
rect 49568 39380 49574 39432
rect 49881 39423 49939 39429
rect 49881 39389 49893 39423
rect 49927 39420 49939 39423
rect 49927 39392 50108 39420
rect 49927 39389 49939 39392
rect 49881 39383 49939 39389
rect 47029 39355 47087 39361
rect 30760 39324 31524 39352
rect 29362 39284 29368 39296
rect 28644 39256 29368 39284
rect 21269 39247 21327 39253
rect 29362 39244 29368 39256
rect 29420 39244 29426 39296
rect 29454 39244 29460 39296
rect 29512 39284 29518 39296
rect 31386 39284 31392 39296
rect 29512 39256 31392 39284
rect 29512 39244 29518 39256
rect 31386 39244 31392 39256
rect 31444 39244 31450 39296
rect 31496 39284 31524 39324
rect 38304 39324 38884 39352
rect 40052 39324 43208 39352
rect 32674 39284 32680 39296
rect 31496 39256 32680 39284
rect 32674 39244 32680 39256
rect 32732 39244 32738 39296
rect 32766 39244 32772 39296
rect 32824 39284 32830 39296
rect 33689 39287 33747 39293
rect 33689 39284 33701 39287
rect 32824 39256 33701 39284
rect 32824 39244 32830 39256
rect 33689 39253 33701 39256
rect 33735 39284 33747 39287
rect 34330 39284 34336 39296
rect 33735 39256 34336 39284
rect 33735 39253 33747 39256
rect 33689 39247 33747 39253
rect 34330 39244 34336 39256
rect 34388 39284 34394 39296
rect 35066 39284 35072 39296
rect 34388 39256 35072 39284
rect 34388 39244 34394 39256
rect 35066 39244 35072 39256
rect 35124 39244 35130 39296
rect 35434 39244 35440 39296
rect 35492 39244 35498 39296
rect 37366 39244 37372 39296
rect 37424 39284 37430 39296
rect 38304 39284 38332 39324
rect 37424 39256 38332 39284
rect 38856 39284 38884 39324
rect 40126 39284 40132 39296
rect 38856 39256 40132 39284
rect 37424 39244 37430 39256
rect 40126 39244 40132 39256
rect 40184 39244 40190 39296
rect 40221 39287 40279 39293
rect 40221 39253 40233 39287
rect 40267 39284 40279 39287
rect 40586 39284 40592 39296
rect 40267 39256 40592 39284
rect 40267 39253 40279 39256
rect 40221 39247 40279 39253
rect 40586 39244 40592 39256
rect 40644 39244 40650 39296
rect 41046 39244 41052 39296
rect 41104 39244 41110 39296
rect 41782 39244 41788 39296
rect 41840 39284 41846 39296
rect 42426 39284 42432 39296
rect 41840 39256 42432 39284
rect 41840 39244 41846 39256
rect 42426 39244 42432 39256
rect 42484 39244 42490 39296
rect 42610 39244 42616 39296
rect 42668 39244 42674 39296
rect 43180 39284 43208 39324
rect 44376 39324 45048 39352
rect 44376 39284 44404 39324
rect 43180 39256 44404 39284
rect 44818 39244 44824 39296
rect 44876 39244 44882 39296
rect 45020 39284 45048 39324
rect 47029 39321 47041 39355
rect 47075 39321 47087 39355
rect 50080 39352 50108 39392
rect 50154 39380 50160 39432
rect 50212 39380 50218 39432
rect 50433 39423 50491 39429
rect 50433 39389 50445 39423
rect 50479 39420 50491 39423
rect 50522 39420 50528 39432
rect 50479 39392 50528 39420
rect 50479 39389 50491 39392
rect 50433 39383 50491 39389
rect 50522 39380 50528 39392
rect 50580 39380 50586 39432
rect 51644 39429 51672 39460
rect 52181 39457 52193 39491
rect 52227 39488 52239 39491
rect 52546 39488 52552 39500
rect 52227 39460 52552 39488
rect 52227 39457 52239 39460
rect 52181 39451 52239 39457
rect 52546 39448 52552 39460
rect 52604 39488 52610 39500
rect 53650 39488 53656 39500
rect 52604 39460 53656 39488
rect 52604 39448 52610 39460
rect 53650 39448 53656 39460
rect 53708 39448 53714 39500
rect 54389 39491 54447 39497
rect 54389 39457 54401 39491
rect 54435 39488 54447 39491
rect 55677 39491 55735 39497
rect 55677 39488 55689 39491
rect 54435 39460 55689 39488
rect 54435 39457 54447 39460
rect 54389 39451 54447 39457
rect 55677 39457 55689 39460
rect 55723 39457 55735 39491
rect 55677 39451 55735 39457
rect 51629 39423 51687 39429
rect 51629 39389 51641 39423
rect 51675 39389 51687 39423
rect 51629 39383 51687 39389
rect 54478 39380 54484 39432
rect 54536 39380 54542 39432
rect 54570 39380 54576 39432
rect 54628 39380 54634 39432
rect 54846 39380 54852 39432
rect 54904 39420 54910 39432
rect 55030 39420 55036 39432
rect 54904 39392 55036 39420
rect 54904 39380 54910 39392
rect 55030 39380 55036 39392
rect 55088 39420 55094 39432
rect 55401 39423 55459 39429
rect 55401 39420 55413 39423
rect 55088 39392 55413 39420
rect 55088 39380 55094 39392
rect 55401 39389 55413 39392
rect 55447 39389 55459 39423
rect 55401 39383 55459 39389
rect 56229 39423 56287 39429
rect 56229 39389 56241 39423
rect 56275 39389 56287 39423
rect 56229 39383 56287 39389
rect 51077 39355 51135 39361
rect 51077 39352 51089 39355
rect 47029 39315 47087 39321
rect 47136 39324 48544 39352
rect 50080 39324 51089 39352
rect 47136 39284 47164 39324
rect 45020 39256 47164 39284
rect 48516 39284 48544 39324
rect 51077 39321 51089 39324
rect 51123 39321 51135 39355
rect 51077 39315 51135 39321
rect 52656 39324 54156 39352
rect 52656 39284 52684 39324
rect 48516 39256 52684 39284
rect 52730 39244 52736 39296
rect 52788 39284 52794 39296
rect 54021 39287 54079 39293
rect 54021 39284 54033 39287
rect 52788 39256 54033 39284
rect 52788 39244 52794 39256
rect 54021 39253 54033 39256
rect 54067 39253 54079 39287
rect 54128 39284 54156 39324
rect 54202 39312 54208 39364
rect 54260 39352 54266 39364
rect 56244 39352 56272 39383
rect 57146 39380 57152 39432
rect 57204 39380 57210 39432
rect 57330 39380 57336 39432
rect 57388 39380 57394 39432
rect 57698 39380 57704 39432
rect 57756 39420 57762 39432
rect 59262 39420 59268 39432
rect 57756 39392 59268 39420
rect 57756 39380 57762 39392
rect 59262 39380 59268 39392
rect 59320 39420 59326 39432
rect 59357 39423 59415 39429
rect 59357 39420 59369 39423
rect 59320 39392 59369 39420
rect 59320 39380 59326 39392
rect 59357 39389 59369 39392
rect 59403 39389 59415 39423
rect 59357 39383 59415 39389
rect 60001 39423 60059 39429
rect 60001 39389 60013 39423
rect 60047 39389 60059 39423
rect 60001 39383 60059 39389
rect 54260 39324 56272 39352
rect 54260 39312 54266 39324
rect 55214 39284 55220 39296
rect 54128 39256 55220 39284
rect 54021 39247 54079 39253
rect 55214 39244 55220 39256
rect 55272 39244 55278 39296
rect 56134 39244 56140 39296
rect 56192 39284 56198 39296
rect 56505 39287 56563 39293
rect 56505 39284 56517 39287
rect 56192 39256 56517 39284
rect 56192 39244 56198 39256
rect 56505 39253 56517 39256
rect 56551 39253 56563 39287
rect 57348 39284 57376 39380
rect 58802 39312 58808 39364
rect 58860 39352 58866 39364
rect 60016 39352 60044 39383
rect 58860 39324 60044 39352
rect 58860 39312 58866 39324
rect 57790 39284 57796 39296
rect 57348 39256 57796 39284
rect 56505 39247 56563 39253
rect 57790 39244 57796 39256
rect 57848 39244 57854 39296
rect 552 39194 66424 39216
rect 552 39142 1998 39194
rect 2050 39142 2062 39194
rect 2114 39142 2126 39194
rect 2178 39142 2190 39194
rect 2242 39142 2254 39194
rect 2306 39142 50998 39194
rect 51050 39142 51062 39194
rect 51114 39142 51126 39194
rect 51178 39142 51190 39194
rect 51242 39142 51254 39194
rect 51306 39142 66424 39194
rect 552 39120 66424 39142
rect 8202 39040 8208 39092
rect 8260 39040 8266 39092
rect 12526 39040 12532 39092
rect 12584 39080 12590 39092
rect 12621 39083 12679 39089
rect 12621 39080 12633 39083
rect 12584 39052 12633 39080
rect 12584 39040 12590 39052
rect 12621 39049 12633 39052
rect 12667 39049 12679 39083
rect 13814 39080 13820 39092
rect 12621 39043 12679 39049
rect 12820 39052 13820 39080
rect 12250 38972 12256 39024
rect 12308 39012 12314 39024
rect 12820 39012 12848 39052
rect 13814 39040 13820 39052
rect 13872 39040 13878 39092
rect 13906 39040 13912 39092
rect 13964 39080 13970 39092
rect 13964 39052 16252 39080
rect 13964 39040 13970 39052
rect 13998 39012 14004 39024
rect 12308 38984 12848 39012
rect 13096 38984 14004 39012
rect 12308 38972 12314 38984
rect 6457 38947 6515 38953
rect 6457 38913 6469 38947
rect 6503 38944 6515 38947
rect 7098 38944 7104 38956
rect 6503 38916 7104 38944
rect 6503 38913 6515 38916
rect 6457 38907 6515 38913
rect 7098 38904 7104 38916
rect 7156 38944 7162 38956
rect 7926 38944 7932 38956
rect 7156 38916 7932 38944
rect 7156 38904 7162 38916
rect 7926 38904 7932 38916
rect 7984 38904 7990 38956
rect 8386 38904 8392 38956
rect 8444 38944 8450 38956
rect 9306 38944 9312 38956
rect 8444 38916 9312 38944
rect 8444 38904 8450 38916
rect 9306 38904 9312 38916
rect 9364 38944 9370 38956
rect 9401 38947 9459 38953
rect 9401 38944 9413 38947
rect 9364 38916 9413 38944
rect 9364 38904 9370 38916
rect 9401 38913 9413 38916
rect 9447 38913 9459 38947
rect 9401 38907 9459 38913
rect 10318 38904 10324 38956
rect 10376 38904 10382 38956
rect 13096 38953 13124 38984
rect 13998 38972 14004 38984
rect 14056 38972 14062 39024
rect 13081 38947 13139 38953
rect 13081 38913 13093 38947
rect 13127 38913 13139 38947
rect 13081 38907 13139 38913
rect 13170 38904 13176 38956
rect 13228 38944 13234 38956
rect 14461 38947 14519 38953
rect 14461 38944 14473 38947
rect 13228 38916 14473 38944
rect 13228 38904 13234 38916
rect 14461 38913 14473 38916
rect 14507 38913 14519 38947
rect 14461 38907 14519 38913
rect 15102 38904 15108 38956
rect 15160 38944 15166 38956
rect 15289 38947 15347 38953
rect 15289 38944 15301 38947
rect 15160 38916 15301 38944
rect 15160 38904 15166 38916
rect 15289 38913 15301 38916
rect 15335 38913 15347 38947
rect 15289 38907 15347 38913
rect 15378 38904 15384 38956
rect 15436 38904 15442 38956
rect 16224 38953 16252 39052
rect 17494 39040 17500 39092
rect 17552 39080 17558 39092
rect 18693 39083 18751 39089
rect 18693 39080 18705 39083
rect 17552 39052 18705 39080
rect 17552 39040 17558 39052
rect 18693 39049 18705 39052
rect 18739 39049 18751 39083
rect 18693 39043 18751 39049
rect 19334 39040 19340 39092
rect 19392 39080 19398 39092
rect 19429 39083 19487 39089
rect 19429 39080 19441 39083
rect 19392 39052 19441 39080
rect 19392 39040 19398 39052
rect 19429 39049 19441 39052
rect 19475 39049 19487 39083
rect 19429 39043 19487 39049
rect 19702 39040 19708 39092
rect 19760 39080 19766 39092
rect 28948 39080 28954 39092
rect 19760 39052 28954 39080
rect 19760 39040 19766 39052
rect 28948 39040 28954 39052
rect 29006 39040 29012 39092
rect 29270 39089 29276 39092
rect 29260 39083 29276 39089
rect 29260 39049 29272 39083
rect 29260 39043 29276 39049
rect 29270 39040 29276 39043
rect 29328 39040 29334 39092
rect 29638 39040 29644 39092
rect 29696 39080 29702 39092
rect 41782 39080 41788 39092
rect 29696 39052 41788 39080
rect 29696 39040 29702 39052
rect 41782 39040 41788 39052
rect 41840 39040 41846 39092
rect 41984 39052 43208 39080
rect 18506 38972 18512 39024
rect 18564 39012 18570 39024
rect 24118 39012 24124 39024
rect 18564 38984 24124 39012
rect 18564 38972 18570 38984
rect 24118 38972 24124 38984
rect 24176 38972 24182 39024
rect 24670 38972 24676 39024
rect 24728 38972 24734 39024
rect 24946 38972 24952 39024
rect 25004 39012 25010 39024
rect 25004 38984 26832 39012
rect 25004 38972 25010 38984
rect 16209 38947 16267 38953
rect 16209 38913 16221 38947
rect 16255 38913 16267 38947
rect 16209 38907 16267 38913
rect 19886 38904 19892 38956
rect 19944 38904 19950 38956
rect 19978 38904 19984 38956
rect 20036 38904 20042 38956
rect 20622 38904 20628 38956
rect 20680 38944 20686 38956
rect 20717 38947 20775 38953
rect 20717 38944 20729 38947
rect 20680 38916 20729 38944
rect 20680 38904 20686 38916
rect 20717 38913 20729 38916
rect 20763 38913 20775 38947
rect 20717 38907 20775 38913
rect 20809 38947 20867 38953
rect 20809 38913 20821 38947
rect 20855 38913 20867 38947
rect 20809 38907 20867 38913
rect 9674 38876 9680 38888
rect 7866 38848 9680 38876
rect 9674 38836 9680 38848
rect 9732 38876 9738 38888
rect 9950 38876 9956 38888
rect 9732 38848 9956 38876
rect 9732 38836 9738 38848
rect 9950 38836 9956 38848
rect 10008 38836 10014 38888
rect 10045 38879 10103 38885
rect 10045 38845 10057 38879
rect 10091 38845 10103 38879
rect 10045 38839 10103 38845
rect 14277 38879 14335 38885
rect 14277 38845 14289 38879
rect 14323 38876 14335 38879
rect 15562 38876 15568 38888
rect 14323 38848 15568 38876
rect 14323 38845 14335 38848
rect 14277 38839 14335 38845
rect 6733 38811 6791 38817
rect 6733 38777 6745 38811
rect 6779 38777 6791 38811
rect 6733 38771 6791 38777
rect 9217 38811 9275 38817
rect 9217 38777 9229 38811
rect 9263 38808 9275 38811
rect 10060 38808 10088 38839
rect 15562 38836 15568 38848
rect 15620 38836 15626 38888
rect 19337 38879 19395 38885
rect 19337 38845 19349 38879
rect 19383 38876 19395 38879
rect 19426 38876 19432 38888
rect 19383 38848 19432 38876
rect 19383 38845 19395 38848
rect 19337 38839 19395 38845
rect 19426 38836 19432 38848
rect 19484 38836 19490 38888
rect 19610 38836 19616 38888
rect 19668 38876 19674 38888
rect 19797 38879 19855 38885
rect 19797 38876 19809 38879
rect 19668 38848 19809 38876
rect 19668 38836 19674 38848
rect 19797 38845 19809 38848
rect 19843 38845 19855 38879
rect 19996 38876 20024 38904
rect 20824 38876 20852 38907
rect 21358 38904 21364 38956
rect 21416 38944 21422 38956
rect 21637 38947 21695 38953
rect 21637 38944 21649 38947
rect 21416 38916 21649 38944
rect 21416 38904 21422 38916
rect 21637 38913 21649 38916
rect 21683 38944 21695 38947
rect 24486 38944 24492 38956
rect 21683 38916 24492 38944
rect 21683 38913 21695 38916
rect 21637 38907 21695 38913
rect 24486 38904 24492 38916
rect 24544 38904 24550 38956
rect 25130 38904 25136 38956
rect 25188 38904 25194 38956
rect 25317 38947 25375 38953
rect 25317 38913 25329 38947
rect 25363 38944 25375 38947
rect 26234 38944 26240 38956
rect 25363 38916 26240 38944
rect 25363 38913 25375 38916
rect 25317 38907 25375 38913
rect 26234 38904 26240 38916
rect 26292 38904 26298 38956
rect 26804 38944 26832 38984
rect 26878 38972 26884 39024
rect 26936 38972 26942 39024
rect 30834 38972 30840 39024
rect 30892 39012 30898 39024
rect 31665 39015 31723 39021
rect 31665 39012 31677 39015
rect 30892 38984 31677 39012
rect 30892 38972 30898 38984
rect 31665 38981 31677 38984
rect 31711 38981 31723 39015
rect 31665 38975 31723 38981
rect 32214 38972 32220 39024
rect 32272 39012 32278 39024
rect 32401 39015 32459 39021
rect 32401 39012 32413 39015
rect 32272 38984 32413 39012
rect 32272 38972 32278 38984
rect 32401 38981 32413 38984
rect 32447 38981 32459 39015
rect 33686 39012 33692 39024
rect 32401 38975 32459 38981
rect 32508 38984 33692 39012
rect 28902 38944 28908 38956
rect 26804 38916 28908 38944
rect 28902 38904 28908 38916
rect 28960 38904 28966 38956
rect 28997 38947 29055 38953
rect 28997 38913 29009 38947
rect 29043 38944 29055 38947
rect 30006 38944 30012 38956
rect 29043 38916 30012 38944
rect 29043 38913 29055 38916
rect 28997 38907 29055 38913
rect 30006 38904 30012 38916
rect 30064 38904 30070 38956
rect 30558 38904 30564 38956
rect 30616 38944 30622 38956
rect 30745 38947 30803 38953
rect 30745 38944 30757 38947
rect 30616 38916 30757 38944
rect 30616 38904 30622 38916
rect 30745 38913 30757 38916
rect 30791 38944 30803 38947
rect 31110 38944 31116 38956
rect 30791 38916 31116 38944
rect 30791 38913 30803 38916
rect 30745 38907 30803 38913
rect 31110 38904 31116 38916
rect 31168 38904 31174 38956
rect 31481 38947 31539 38953
rect 31481 38913 31493 38947
rect 31527 38944 31539 38947
rect 32122 38944 32128 38956
rect 31527 38916 32128 38944
rect 31527 38913 31539 38916
rect 31481 38907 31539 38913
rect 32122 38904 32128 38916
rect 32180 38904 32186 38956
rect 32508 38944 32536 38984
rect 33686 38972 33692 38984
rect 33744 38972 33750 39024
rect 34054 38972 34060 39024
rect 34112 39012 34118 39024
rect 34149 39015 34207 39021
rect 34149 39012 34161 39015
rect 34112 38984 34161 39012
rect 34112 38972 34118 38984
rect 34149 38981 34161 38984
rect 34195 39012 34207 39015
rect 34606 39012 34612 39024
rect 34195 38984 34612 39012
rect 34195 38981 34207 38984
rect 34149 38975 34207 38981
rect 34606 38972 34612 38984
rect 34664 38972 34670 39024
rect 39114 39012 39120 39024
rect 37292 38984 39120 39012
rect 32232 38916 32536 38944
rect 33045 38947 33103 38953
rect 19996 38848 20852 38876
rect 19797 38839 19855 38845
rect 21082 38836 21088 38888
rect 21140 38876 21146 38888
rect 21453 38879 21511 38885
rect 21453 38876 21465 38879
rect 21140 38848 21465 38876
rect 21140 38836 21146 38848
rect 21453 38845 21465 38848
rect 21499 38876 21511 38879
rect 22465 38879 22523 38885
rect 22465 38876 22477 38879
rect 21499 38848 22477 38876
rect 21499 38845 21511 38848
rect 21453 38839 21511 38845
rect 22465 38845 22477 38848
rect 22511 38845 22523 38879
rect 22465 38839 22523 38845
rect 23474 38836 23480 38888
rect 23532 38876 23538 38888
rect 23569 38879 23627 38885
rect 23569 38876 23581 38879
rect 23532 38848 23581 38876
rect 23532 38836 23538 38848
rect 23569 38845 23581 38848
rect 23615 38876 23627 38879
rect 24213 38879 24271 38885
rect 24213 38876 24225 38879
rect 23615 38848 24225 38876
rect 23615 38845 23627 38848
rect 23569 38839 23627 38845
rect 24213 38845 24225 38848
rect 24259 38845 24271 38879
rect 24213 38839 24271 38845
rect 25038 38836 25044 38888
rect 25096 38836 25102 38888
rect 25501 38879 25559 38885
rect 25501 38876 25513 38879
rect 25332 38848 25513 38876
rect 10226 38808 10232 38820
rect 9263 38780 9996 38808
rect 10060 38780 10232 38808
rect 9263 38777 9275 38780
rect 9217 38771 9275 38777
rect 6748 38740 6776 38771
rect 6914 38740 6920 38752
rect 6748 38712 6920 38740
rect 6914 38700 6920 38712
rect 6972 38700 6978 38752
rect 7006 38700 7012 38752
rect 7064 38740 7070 38752
rect 8849 38743 8907 38749
rect 8849 38740 8861 38743
rect 7064 38712 8861 38740
rect 7064 38700 7070 38712
rect 8849 38709 8861 38712
rect 8895 38709 8907 38743
rect 8849 38703 8907 38709
rect 9309 38743 9367 38749
rect 9309 38709 9321 38743
rect 9355 38740 9367 38743
rect 9858 38740 9864 38752
rect 9355 38712 9864 38740
rect 9355 38709 9367 38712
rect 9309 38703 9367 38709
rect 9858 38700 9864 38712
rect 9916 38700 9922 38752
rect 9968 38740 9996 38780
rect 10226 38768 10232 38780
rect 10284 38768 10290 38820
rect 10318 38768 10324 38820
rect 10376 38808 10382 38820
rect 10376 38780 10810 38808
rect 10376 38768 10382 38780
rect 12066 38768 12072 38820
rect 12124 38768 12130 38820
rect 12989 38811 13047 38817
rect 12989 38777 13001 38811
rect 13035 38808 13047 38811
rect 15657 38811 15715 38817
rect 15657 38808 15669 38811
rect 13035 38780 15669 38808
rect 13035 38777 13047 38780
rect 12989 38771 13047 38777
rect 15657 38777 15669 38780
rect 15703 38777 15715 38811
rect 15657 38771 15715 38777
rect 16206 38768 16212 38820
rect 16264 38808 16270 38820
rect 16761 38811 16819 38817
rect 16761 38808 16773 38811
rect 16264 38780 16773 38808
rect 16264 38768 16270 38780
rect 16761 38777 16773 38780
rect 16807 38777 16819 38811
rect 16761 38771 16819 38777
rect 18509 38811 18567 38817
rect 18509 38777 18521 38811
rect 18555 38808 18567 38811
rect 20530 38808 20536 38820
rect 18555 38780 20536 38808
rect 18555 38777 18567 38780
rect 18509 38771 18567 38777
rect 20530 38768 20536 38780
rect 20588 38768 20594 38820
rect 20625 38811 20683 38817
rect 20625 38777 20637 38811
rect 20671 38808 20683 38811
rect 21913 38811 21971 38817
rect 21913 38808 21925 38811
rect 20671 38780 21925 38808
rect 20671 38777 20683 38780
rect 20625 38771 20683 38777
rect 21913 38777 21925 38780
rect 21959 38777 21971 38811
rect 21913 38771 21971 38777
rect 23198 38768 23204 38820
rect 23256 38808 23262 38820
rect 24305 38811 24363 38817
rect 23256 38780 23980 38808
rect 23256 38768 23262 38780
rect 10962 38740 10968 38752
rect 9968 38712 10968 38740
rect 10962 38700 10968 38712
rect 11020 38700 11026 38752
rect 13814 38700 13820 38752
rect 13872 38740 13878 38752
rect 13909 38743 13967 38749
rect 13909 38740 13921 38743
rect 13872 38712 13921 38740
rect 13872 38700 13878 38712
rect 13909 38709 13921 38712
rect 13955 38709 13967 38743
rect 13909 38703 13967 38709
rect 14369 38743 14427 38749
rect 14369 38709 14381 38743
rect 14415 38740 14427 38743
rect 14829 38743 14887 38749
rect 14829 38740 14841 38743
rect 14415 38712 14841 38740
rect 14415 38709 14427 38712
rect 14369 38703 14427 38709
rect 14829 38709 14841 38712
rect 14875 38709 14887 38743
rect 14829 38703 14887 38709
rect 15197 38743 15255 38749
rect 15197 38709 15209 38743
rect 15243 38740 15255 38743
rect 15378 38740 15384 38752
rect 15243 38712 15384 38740
rect 15243 38709 15255 38712
rect 15197 38703 15255 38709
rect 15378 38700 15384 38712
rect 15436 38740 15442 38752
rect 16390 38740 16396 38752
rect 15436 38712 16396 38740
rect 15436 38700 15442 38712
rect 16390 38700 16396 38712
rect 16448 38700 16454 38752
rect 20254 38700 20260 38752
rect 20312 38700 20318 38752
rect 20346 38700 20352 38752
rect 20404 38740 20410 38752
rect 20714 38740 20720 38752
rect 20404 38712 20720 38740
rect 20404 38700 20410 38712
rect 20714 38700 20720 38712
rect 20772 38700 20778 38752
rect 20806 38700 20812 38752
rect 20864 38740 20870 38752
rect 21085 38743 21143 38749
rect 21085 38740 21097 38743
rect 20864 38712 21097 38740
rect 20864 38700 20870 38712
rect 21085 38709 21097 38712
rect 21131 38709 21143 38743
rect 21085 38703 21143 38709
rect 21545 38743 21603 38749
rect 21545 38709 21557 38743
rect 21591 38740 21603 38743
rect 21818 38740 21824 38752
rect 21591 38712 21824 38740
rect 21591 38709 21603 38712
rect 21545 38703 21603 38709
rect 21818 38700 21824 38712
rect 21876 38700 21882 38752
rect 23014 38700 23020 38752
rect 23072 38700 23078 38752
rect 23750 38700 23756 38752
rect 23808 38740 23814 38752
rect 23845 38743 23903 38749
rect 23845 38740 23857 38743
rect 23808 38712 23857 38740
rect 23808 38700 23814 38712
rect 23845 38709 23857 38712
rect 23891 38709 23903 38743
rect 23952 38740 23980 38780
rect 24305 38777 24317 38811
rect 24351 38808 24363 38811
rect 25332 38808 25360 38848
rect 25501 38845 25513 38848
rect 25547 38845 25559 38879
rect 25501 38839 25559 38845
rect 26142 38836 26148 38888
rect 26200 38836 26206 38888
rect 26329 38879 26387 38885
rect 26329 38845 26341 38879
rect 26375 38876 26387 38879
rect 27614 38876 27620 38888
rect 26375 38848 27620 38876
rect 26375 38845 26387 38848
rect 26329 38839 26387 38845
rect 27614 38836 27620 38848
rect 27672 38876 27678 38888
rect 28534 38876 28540 38888
rect 27672 38848 28540 38876
rect 27672 38836 27678 38848
rect 28534 38836 28540 38848
rect 28592 38836 28598 38888
rect 32232 38876 32260 38916
rect 33045 38913 33057 38947
rect 33091 38944 33103 38947
rect 33962 38944 33968 38956
rect 33091 38916 33968 38944
rect 33091 38913 33103 38916
rect 33045 38907 33103 38913
rect 30760 38848 32260 38876
rect 32309 38879 32367 38885
rect 27798 38808 27804 38820
rect 24351 38780 25360 38808
rect 25608 38780 27804 38808
rect 24351 38777 24363 38780
rect 24305 38771 24363 38777
rect 25608 38740 25636 38780
rect 27798 38768 27804 38780
rect 27856 38768 27862 38820
rect 28626 38768 28632 38820
rect 28684 38808 28690 38820
rect 28684 38780 29762 38808
rect 28684 38768 28690 38780
rect 23952 38712 25636 38740
rect 23845 38703 23903 38709
rect 25682 38700 25688 38752
rect 25740 38740 25746 38752
rect 28948 38740 28954 38752
rect 25740 38712 28954 38740
rect 25740 38700 25746 38712
rect 28948 38700 28954 38712
rect 29006 38700 29012 38752
rect 29086 38700 29092 38752
rect 29144 38740 29150 38752
rect 30760 38740 30788 38848
rect 32309 38845 32321 38879
rect 32355 38876 32367 38879
rect 32861 38879 32919 38885
rect 32861 38876 32873 38879
rect 32355 38848 32873 38876
rect 32355 38845 32367 38848
rect 32309 38839 32367 38845
rect 32861 38845 32873 38848
rect 32907 38845 32919 38879
rect 32861 38839 32919 38845
rect 31570 38808 31576 38820
rect 31220 38780 31576 38808
rect 31220 38752 31248 38780
rect 31570 38768 31576 38780
rect 31628 38808 31634 38820
rect 32324 38808 32352 38839
rect 31628 38780 32352 38808
rect 31628 38768 31634 38780
rect 32766 38768 32772 38820
rect 32824 38768 32830 38820
rect 29144 38712 30788 38740
rect 29144 38700 29150 38712
rect 30834 38700 30840 38752
rect 30892 38700 30898 38752
rect 31202 38700 31208 38752
rect 31260 38700 31266 38752
rect 31297 38743 31355 38749
rect 31297 38709 31309 38743
rect 31343 38740 31355 38743
rect 31386 38740 31392 38752
rect 31343 38712 31392 38740
rect 31343 38709 31355 38712
rect 31297 38703 31355 38709
rect 31386 38700 31392 38712
rect 31444 38700 31450 38752
rect 32122 38700 32128 38752
rect 32180 38740 32186 38752
rect 33060 38740 33088 38907
rect 33962 38904 33968 38916
rect 34020 38904 34026 38956
rect 35897 38947 35955 38953
rect 35897 38913 35909 38947
rect 35943 38944 35955 38947
rect 37182 38944 37188 38956
rect 35943 38916 37188 38944
rect 35943 38913 35955 38916
rect 35897 38907 35955 38913
rect 37182 38904 37188 38916
rect 37240 38904 37246 38956
rect 37292 38953 37320 38984
rect 39114 38972 39120 38984
rect 39172 38972 39178 39024
rect 39298 38972 39304 39024
rect 39356 38972 39362 39024
rect 40126 38972 40132 39024
rect 40184 39012 40190 39024
rect 40184 38984 40724 39012
rect 40184 38972 40190 38984
rect 37277 38947 37335 38953
rect 37277 38913 37289 38947
rect 37323 38913 37335 38947
rect 37277 38907 37335 38913
rect 37366 38904 37372 38956
rect 37424 38904 37430 38956
rect 38194 38944 38200 38956
rect 37476 38916 38200 38944
rect 37476 38876 37504 38916
rect 38194 38904 38200 38916
rect 38252 38904 38258 38956
rect 38286 38904 38292 38956
rect 38344 38904 38350 38956
rect 38470 38904 38476 38956
rect 38528 38944 38534 38956
rect 39025 38947 39083 38953
rect 39025 38944 39037 38947
rect 38528 38916 39037 38944
rect 38528 38904 38534 38916
rect 39025 38913 39037 38916
rect 39071 38913 39083 38947
rect 39025 38907 39083 38913
rect 39945 38947 40003 38953
rect 39945 38913 39957 38947
rect 39991 38944 40003 38947
rect 40218 38944 40224 38956
rect 39991 38916 40224 38944
rect 39991 38913 40003 38916
rect 39945 38907 40003 38913
rect 40218 38904 40224 38916
rect 40276 38904 40282 38956
rect 40586 38904 40592 38956
rect 40644 38904 40650 38956
rect 40696 38953 40724 38984
rect 40681 38947 40739 38953
rect 40681 38913 40693 38947
rect 40727 38944 40739 38947
rect 41230 38944 41236 38956
rect 40727 38916 41236 38944
rect 40727 38913 40739 38916
rect 40681 38907 40739 38913
rect 41230 38904 41236 38916
rect 41288 38944 41294 38956
rect 41984 38944 42012 39052
rect 41288 38916 42012 38944
rect 41288 38904 41294 38916
rect 42886 38904 42892 38956
rect 42944 38944 42950 38956
rect 42981 38947 43039 38953
rect 42981 38944 42993 38947
rect 42944 38916 42993 38944
rect 42944 38904 42950 38916
rect 42981 38913 42993 38916
rect 43027 38913 43039 38947
rect 43180 38944 43208 39052
rect 43438 39040 43444 39092
rect 43496 39080 43502 39092
rect 43533 39083 43591 39089
rect 43533 39080 43545 39083
rect 43496 39052 43545 39080
rect 43496 39040 43502 39052
rect 43533 39049 43545 39052
rect 43579 39049 43591 39083
rect 43533 39043 43591 39049
rect 45833 39083 45891 39089
rect 45833 39049 45845 39083
rect 45879 39080 45891 39083
rect 47486 39080 47492 39092
rect 45879 39052 47492 39080
rect 45879 39049 45891 39052
rect 45833 39043 45891 39049
rect 47486 39040 47492 39052
rect 47544 39040 47550 39092
rect 47670 39040 47676 39092
rect 47728 39080 47734 39092
rect 48314 39080 48320 39092
rect 47728 39052 48320 39080
rect 47728 39040 47734 39052
rect 48314 39040 48320 39052
rect 48372 39040 48378 39092
rect 48958 39040 48964 39092
rect 49016 39080 49022 39092
rect 50433 39083 50491 39089
rect 50433 39080 50445 39083
rect 49016 39052 50445 39080
rect 49016 39040 49022 39052
rect 50433 39049 50445 39052
rect 50479 39049 50491 39083
rect 50433 39043 50491 39049
rect 54202 39040 54208 39092
rect 54260 39040 54266 39092
rect 54478 39040 54484 39092
rect 54536 39080 54542 39092
rect 54757 39083 54815 39089
rect 54757 39080 54769 39083
rect 54536 39052 54769 39080
rect 54536 39040 54542 39052
rect 54757 39049 54769 39052
rect 54803 39049 54815 39083
rect 57320 39083 57378 39089
rect 54757 39043 54815 39049
rect 55140 39052 56272 39080
rect 43622 38972 43628 39024
rect 43680 39012 43686 39024
rect 50338 39012 50344 39024
rect 43680 38984 46060 39012
rect 43680 38972 43686 38984
rect 43990 38944 43996 38956
rect 43180 38916 43996 38944
rect 42981 38907 43039 38913
rect 43990 38904 43996 38916
rect 44048 38944 44054 38956
rect 44085 38947 44143 38953
rect 44085 38944 44097 38947
rect 44048 38916 44097 38944
rect 44048 38904 44054 38916
rect 44085 38913 44097 38916
rect 44131 38913 44143 38947
rect 44085 38907 44143 38913
rect 45189 38947 45247 38953
rect 45189 38913 45201 38947
rect 45235 38944 45247 38947
rect 45554 38944 45560 38956
rect 45235 38916 45560 38944
rect 45235 38913 45247 38916
rect 45189 38907 45247 38913
rect 45554 38904 45560 38916
rect 45612 38904 45618 38956
rect 45925 38947 45983 38953
rect 45925 38944 45937 38947
rect 45664 38916 45937 38944
rect 35912 38848 37504 38876
rect 38013 38879 38071 38885
rect 33962 38768 33968 38820
rect 34020 38808 34026 38820
rect 34146 38808 34152 38820
rect 34020 38780 34152 38808
rect 34020 38768 34026 38780
rect 34146 38768 34152 38780
rect 34204 38808 34210 38820
rect 34204 38780 34454 38808
rect 34204 38768 34210 38780
rect 35618 38768 35624 38820
rect 35676 38768 35682 38820
rect 32180 38712 33088 38740
rect 32180 38700 32186 38712
rect 34330 38700 34336 38752
rect 34388 38740 34394 38752
rect 35912 38740 35940 38848
rect 38013 38845 38025 38879
rect 38059 38876 38071 38879
rect 38488 38876 38516 38904
rect 38059 38848 38516 38876
rect 38059 38845 38071 38848
rect 38013 38839 38071 38845
rect 38930 38836 38936 38888
rect 38988 38876 38994 38888
rect 39761 38879 39819 38885
rect 39761 38876 39773 38879
rect 38988 38848 39773 38876
rect 38988 38836 38994 38848
rect 39761 38845 39773 38848
rect 39807 38845 39819 38879
rect 39761 38839 39819 38845
rect 40497 38879 40555 38885
rect 40497 38845 40509 38879
rect 40543 38876 40555 38879
rect 41046 38876 41052 38888
rect 40543 38848 41052 38876
rect 40543 38845 40555 38848
rect 40497 38839 40555 38845
rect 41046 38836 41052 38848
rect 41104 38836 41110 38888
rect 41874 38836 41880 38888
rect 41932 38836 41938 38888
rect 43257 38879 43315 38885
rect 43257 38845 43269 38879
rect 43303 38876 43315 38879
rect 43346 38876 43352 38888
rect 43303 38848 43352 38876
rect 43303 38845 43315 38848
rect 43257 38839 43315 38845
rect 43346 38836 43352 38848
rect 43404 38876 43410 38888
rect 45278 38876 45284 38888
rect 43404 38848 45284 38876
rect 43404 38836 43410 38848
rect 45278 38836 45284 38848
rect 45336 38876 45342 38888
rect 45664 38876 45692 38916
rect 45925 38913 45937 38916
rect 45971 38913 45983 38947
rect 46032 38944 46060 38984
rect 48148 38984 50344 39012
rect 48148 38944 48176 38984
rect 46032 38916 48176 38944
rect 45925 38907 45983 38913
rect 48314 38904 48320 38956
rect 48372 38904 48378 38956
rect 49160 38953 49188 38984
rect 50338 38972 50344 38984
rect 50396 39012 50402 39024
rect 50614 39012 50620 39024
rect 50396 38984 50620 39012
rect 50396 38972 50402 38984
rect 50614 38972 50620 38984
rect 50672 39012 50678 39024
rect 50672 38984 50936 39012
rect 50672 38972 50678 38984
rect 49145 38947 49203 38953
rect 49145 38913 49157 38947
rect 49191 38913 49203 38947
rect 49145 38907 49203 38913
rect 49326 38904 49332 38956
rect 49384 38904 49390 38956
rect 49786 38904 49792 38956
rect 49844 38944 49850 38956
rect 50798 38944 50804 38956
rect 49844 38916 50804 38944
rect 49844 38904 49850 38916
rect 50798 38904 50804 38916
rect 50856 38904 50862 38956
rect 50908 38953 50936 38984
rect 54570 38972 54576 39024
rect 54628 39012 54634 39024
rect 55140 39012 55168 39052
rect 55585 39015 55643 39021
rect 55585 39012 55597 39015
rect 54628 38984 55168 39012
rect 55232 38984 55597 39012
rect 54628 38972 54634 38984
rect 55232 38956 55260 38984
rect 55585 38981 55597 38984
rect 55631 38981 55643 39015
rect 55585 38975 55643 38981
rect 50893 38947 50951 38953
rect 50893 38913 50905 38947
rect 50939 38913 50951 38947
rect 50893 38907 50951 38913
rect 50985 38947 51043 38953
rect 50985 38913 50997 38947
rect 51031 38913 51043 38947
rect 50985 38907 51043 38913
rect 45336 38848 45692 38876
rect 45336 38836 45342 38848
rect 48406 38836 48412 38888
rect 48464 38876 48470 38888
rect 49053 38879 49111 38885
rect 49053 38876 49065 38879
rect 48464 38848 49065 38876
rect 48464 38836 48470 38848
rect 49053 38845 49065 38848
rect 49099 38845 49111 38879
rect 49053 38839 49111 38845
rect 49510 38836 49516 38888
rect 49568 38876 49574 38888
rect 50249 38879 50307 38885
rect 50249 38876 50261 38879
rect 49568 38848 50261 38876
rect 49568 38836 49574 38848
rect 50249 38845 50261 38848
rect 50295 38845 50307 38879
rect 50249 38839 50307 38845
rect 37185 38811 37243 38817
rect 37185 38777 37197 38811
rect 37231 38808 37243 38811
rect 38473 38811 38531 38817
rect 38473 38808 38485 38811
rect 37231 38780 38485 38808
rect 37231 38777 37243 38780
rect 37185 38771 37243 38777
rect 38473 38777 38485 38780
rect 38519 38777 38531 38811
rect 41690 38808 41696 38820
rect 38473 38771 38531 38777
rect 38580 38780 41696 38808
rect 34388 38712 35940 38740
rect 36817 38743 36875 38749
rect 34388 38700 34394 38712
rect 36817 38709 36829 38743
rect 36863 38740 36875 38743
rect 36998 38740 37004 38752
rect 36863 38712 37004 38740
rect 36863 38709 36875 38712
rect 36817 38703 36875 38709
rect 36998 38700 37004 38712
rect 37056 38700 37062 38752
rect 37458 38700 37464 38752
rect 37516 38740 37522 38752
rect 37645 38743 37703 38749
rect 37645 38740 37657 38743
rect 37516 38712 37657 38740
rect 37516 38700 37522 38712
rect 37645 38709 37657 38712
rect 37691 38709 37703 38743
rect 37645 38703 37703 38709
rect 38010 38700 38016 38752
rect 38068 38740 38074 38752
rect 38105 38743 38163 38749
rect 38105 38740 38117 38743
rect 38068 38712 38117 38740
rect 38068 38700 38074 38712
rect 38105 38709 38117 38712
rect 38151 38709 38163 38743
rect 38105 38703 38163 38709
rect 38194 38700 38200 38752
rect 38252 38740 38258 38752
rect 38580 38740 38608 38780
rect 41690 38768 41696 38780
rect 41748 38768 41754 38820
rect 43901 38811 43959 38817
rect 43901 38777 43913 38811
rect 43947 38808 43959 38811
rect 45186 38808 45192 38820
rect 43947 38780 45192 38808
rect 43947 38777 43959 38780
rect 43901 38771 43959 38777
rect 45186 38768 45192 38780
rect 45244 38768 45250 38820
rect 45462 38768 45468 38820
rect 45520 38768 45526 38820
rect 46198 38768 46204 38820
rect 46256 38768 46262 38820
rect 46658 38768 46664 38820
rect 46716 38768 46722 38820
rect 47486 38768 47492 38820
rect 47544 38808 47550 38820
rect 49694 38808 49700 38820
rect 47544 38780 49700 38808
rect 47544 38768 47550 38780
rect 49694 38768 49700 38780
rect 49752 38768 49758 38820
rect 50264 38808 50292 38839
rect 50522 38836 50528 38888
rect 50580 38876 50586 38888
rect 51000 38876 51028 38907
rect 52454 38904 52460 38956
rect 52512 38944 52518 38956
rect 53466 38944 53472 38956
rect 52512 38916 53472 38944
rect 52512 38904 52518 38916
rect 53466 38904 53472 38916
rect 53524 38904 53530 38956
rect 55214 38904 55220 38956
rect 55272 38904 55278 38956
rect 55401 38947 55459 38953
rect 55401 38913 55413 38947
rect 55447 38944 55459 38947
rect 55674 38944 55680 38956
rect 55447 38916 55680 38944
rect 55447 38913 55459 38916
rect 55401 38907 55459 38913
rect 55674 38904 55680 38916
rect 55732 38944 55738 38956
rect 56244 38944 56272 39052
rect 57320 39049 57332 39083
rect 57366 39080 57378 39083
rect 58066 39080 58072 39092
rect 57366 39052 58072 39080
rect 57366 39049 57378 39052
rect 57320 39043 57378 39049
rect 58066 39040 58072 39052
rect 58124 39040 58130 39092
rect 58802 39040 58808 39092
rect 58860 39040 58866 39092
rect 58894 39040 58900 39092
rect 58952 39040 58958 39092
rect 56321 38947 56379 38953
rect 56321 38944 56333 38947
rect 55732 38916 56088 38944
rect 56244 38916 56333 38944
rect 55732 38904 55738 38916
rect 50580 38848 51028 38876
rect 50580 38836 50586 38848
rect 52270 38836 52276 38888
rect 52328 38836 52334 38888
rect 53834 38836 53840 38888
rect 53892 38876 53898 38888
rect 55122 38876 55128 38888
rect 53892 38848 55128 38876
rect 53892 38836 53898 38848
rect 55122 38836 55128 38848
rect 55180 38876 55186 38888
rect 55950 38876 55956 38888
rect 55180 38848 55956 38876
rect 55180 38836 55186 38848
rect 55950 38836 55956 38848
rect 56008 38836 56014 38888
rect 50706 38808 50712 38820
rect 50264 38780 50712 38808
rect 50706 38768 50712 38780
rect 50764 38808 50770 38820
rect 50801 38811 50859 38817
rect 50801 38808 50813 38811
rect 50764 38780 50813 38808
rect 50764 38768 50770 38780
rect 50801 38777 50813 38780
rect 50847 38777 50859 38811
rect 50801 38771 50859 38777
rect 52730 38768 52736 38820
rect 52788 38768 52794 38820
rect 56060 38808 56088 38916
rect 56321 38913 56333 38916
rect 56367 38913 56379 38947
rect 56321 38907 56379 38913
rect 56502 38904 56508 38956
rect 56560 38944 56566 38956
rect 57057 38947 57115 38953
rect 57057 38944 57069 38947
rect 56560 38916 57069 38944
rect 56560 38904 56566 38916
rect 57057 38913 57069 38916
rect 57103 38944 57115 38947
rect 57974 38944 57980 38956
rect 57103 38916 57980 38944
rect 57103 38913 57115 38916
rect 57057 38907 57115 38913
rect 57974 38904 57980 38916
rect 58032 38904 58038 38956
rect 59446 38904 59452 38956
rect 59504 38904 59510 38956
rect 56134 38836 56140 38888
rect 56192 38836 56198 38888
rect 59262 38836 59268 38888
rect 59320 38836 59326 38888
rect 56060 38780 56364 38808
rect 38252 38712 38608 38740
rect 38252 38700 38258 38712
rect 39666 38700 39672 38752
rect 39724 38700 39730 38752
rect 39850 38700 39856 38752
rect 39908 38740 39914 38752
rect 40129 38743 40187 38749
rect 40129 38740 40141 38743
rect 39908 38712 40141 38740
rect 39908 38700 39914 38712
rect 40129 38709 40141 38712
rect 40175 38709 40187 38743
rect 40129 38703 40187 38709
rect 41506 38700 41512 38752
rect 41564 38740 41570 38752
rect 42242 38740 42248 38752
rect 41564 38712 42248 38740
rect 41564 38700 41570 38712
rect 42242 38700 42248 38712
rect 42300 38700 42306 38752
rect 43993 38743 44051 38749
rect 43993 38709 44005 38743
rect 44039 38740 44051 38743
rect 44174 38740 44180 38752
rect 44039 38712 44180 38740
rect 44039 38709 44051 38712
rect 43993 38703 44051 38709
rect 44174 38700 44180 38712
rect 44232 38700 44238 38752
rect 45370 38700 45376 38752
rect 45428 38700 45434 38752
rect 45554 38700 45560 38752
rect 45612 38740 45618 38752
rect 47118 38740 47124 38752
rect 45612 38712 47124 38740
rect 45612 38700 45618 38712
rect 47118 38700 47124 38712
rect 47176 38700 47182 38752
rect 47762 38700 47768 38752
rect 47820 38700 47826 38752
rect 48685 38743 48743 38749
rect 48685 38709 48697 38743
rect 48731 38740 48743 38743
rect 48958 38740 48964 38752
rect 48731 38712 48964 38740
rect 48731 38709 48743 38712
rect 48685 38703 48743 38709
rect 48958 38700 48964 38712
rect 49016 38700 49022 38752
rect 50982 38700 50988 38752
rect 51040 38740 51046 38752
rect 51721 38743 51779 38749
rect 51721 38740 51733 38743
rect 51040 38712 51733 38740
rect 51040 38700 51046 38712
rect 51721 38709 51733 38712
rect 51767 38709 51779 38743
rect 51721 38703 51779 38709
rect 54110 38700 54116 38752
rect 54168 38740 54174 38752
rect 55122 38740 55128 38752
rect 54168 38712 55128 38740
rect 54168 38700 54174 38712
rect 55122 38700 55128 38712
rect 55180 38700 55186 38752
rect 55766 38700 55772 38752
rect 55824 38700 55830 38752
rect 56226 38700 56232 38752
rect 56284 38700 56290 38752
rect 56336 38740 56364 38780
rect 58342 38768 58348 38820
rect 58400 38768 58406 38820
rect 63678 38808 63684 38820
rect 58820 38780 63684 38808
rect 58820 38740 58848 38780
rect 63678 38768 63684 38780
rect 63736 38768 63742 38820
rect 56336 38712 58848 38740
rect 59262 38700 59268 38752
rect 59320 38740 59326 38752
rect 59357 38743 59415 38749
rect 59357 38740 59369 38743
rect 59320 38712 59369 38740
rect 59320 38700 59326 38712
rect 59357 38709 59369 38712
rect 59403 38709 59415 38743
rect 59357 38703 59415 38709
rect 552 38650 66424 38672
rect 552 38598 2918 38650
rect 2970 38598 2982 38650
rect 3034 38598 3046 38650
rect 3098 38598 3110 38650
rect 3162 38598 3174 38650
rect 3226 38598 51918 38650
rect 51970 38598 51982 38650
rect 52034 38598 52046 38650
rect 52098 38598 52110 38650
rect 52162 38598 52174 38650
rect 52226 38598 66424 38650
rect 552 38576 66424 38598
rect 6914 38496 6920 38548
rect 6972 38496 6978 38548
rect 7285 38539 7343 38545
rect 7285 38505 7297 38539
rect 7331 38536 7343 38539
rect 7834 38536 7840 38548
rect 7331 38508 7840 38536
rect 7331 38505 7343 38508
rect 7285 38499 7343 38505
rect 7834 38496 7840 38508
rect 7892 38496 7898 38548
rect 8113 38539 8171 38545
rect 8113 38505 8125 38539
rect 8159 38536 8171 38539
rect 8202 38536 8208 38548
rect 8159 38508 8208 38536
rect 8159 38505 8171 38508
rect 8113 38499 8171 38505
rect 8202 38496 8208 38508
rect 8260 38496 8266 38548
rect 8754 38536 8760 38548
rect 8588 38508 8760 38536
rect 8386 38400 8392 38412
rect 7576 38372 8392 38400
rect 7374 38292 7380 38344
rect 7432 38292 7438 38344
rect 7576 38341 7604 38372
rect 8386 38360 8392 38372
rect 8444 38360 8450 38412
rect 8478 38360 8484 38412
rect 8536 38400 8542 38412
rect 8588 38409 8616 38508
rect 8754 38496 8760 38508
rect 8812 38536 8818 38548
rect 8812 38508 10272 38536
rect 8812 38496 8818 38508
rect 10244 38480 10272 38508
rect 10962 38496 10968 38548
rect 11020 38496 11026 38548
rect 11054 38496 11060 38548
rect 11112 38536 11118 38548
rect 11701 38539 11759 38545
rect 11701 38536 11713 38539
rect 11112 38508 11713 38536
rect 11112 38496 11118 38508
rect 11701 38505 11713 38508
rect 11747 38505 11759 38539
rect 15194 38536 15200 38548
rect 11701 38499 11759 38505
rect 13372 38508 15200 38536
rect 10226 38428 10232 38480
rect 10284 38468 10290 38480
rect 13372 38468 13400 38508
rect 15194 38496 15200 38508
rect 15252 38496 15258 38548
rect 15289 38539 15347 38545
rect 15289 38505 15301 38539
rect 15335 38536 15347 38539
rect 15562 38536 15568 38548
rect 15335 38508 15568 38536
rect 15335 38505 15347 38508
rect 15289 38499 15347 38505
rect 15562 38496 15568 38508
rect 15620 38496 15626 38548
rect 16485 38539 16543 38545
rect 16485 38536 16497 38539
rect 15948 38508 16497 38536
rect 10284 38440 13400 38468
rect 10284 38428 10290 38440
rect 8573 38403 8631 38409
rect 8573 38400 8585 38403
rect 8536 38372 8585 38400
rect 8536 38360 8542 38372
rect 8573 38369 8585 38372
rect 8619 38369 8631 38403
rect 8573 38363 8631 38369
rect 9950 38360 9956 38412
rect 10008 38400 10014 38412
rect 10318 38400 10324 38412
rect 10008 38372 10324 38400
rect 10008 38360 10014 38372
rect 10318 38360 10324 38372
rect 10376 38360 10382 38412
rect 10597 38403 10655 38409
rect 10597 38369 10609 38403
rect 10643 38400 10655 38403
rect 11422 38400 11428 38412
rect 10643 38372 11428 38400
rect 10643 38369 10655 38372
rect 10597 38363 10655 38369
rect 7561 38335 7619 38341
rect 7561 38301 7573 38335
rect 7607 38301 7619 38335
rect 7561 38295 7619 38301
rect 7926 38292 7932 38344
rect 7984 38292 7990 38344
rect 8021 38335 8079 38341
rect 8021 38301 8033 38335
rect 8067 38301 8079 38335
rect 8849 38335 8907 38341
rect 8849 38332 8861 38335
rect 8021 38295 8079 38301
rect 8496 38304 8861 38332
rect 8036 38196 8064 38295
rect 8496 38273 8524 38304
rect 8849 38301 8861 38304
rect 8895 38301 8907 38335
rect 8849 38295 8907 38301
rect 8481 38267 8539 38273
rect 8481 38233 8493 38267
rect 8527 38233 8539 38267
rect 8481 38227 8539 38233
rect 9950 38224 9956 38276
rect 10008 38264 10014 38276
rect 10612 38264 10640 38363
rect 11422 38360 11428 38372
rect 11480 38360 11486 38412
rect 12066 38360 12072 38412
rect 12124 38360 12130 38412
rect 12710 38400 12716 38412
rect 12176 38372 12716 38400
rect 12176 38344 12204 38372
rect 12710 38360 12716 38372
rect 12768 38360 12774 38412
rect 13372 38409 13400 38440
rect 14274 38428 14280 38480
rect 14332 38428 14338 38480
rect 12897 38403 12955 38409
rect 12897 38369 12909 38403
rect 12943 38369 12955 38403
rect 12897 38363 12955 38369
rect 13357 38403 13415 38409
rect 13357 38369 13369 38403
rect 13403 38369 13415 38403
rect 13357 38363 13415 38369
rect 11514 38292 11520 38344
rect 11572 38292 11578 38344
rect 12158 38292 12164 38344
rect 12216 38292 12222 38344
rect 12250 38292 12256 38344
rect 12308 38292 12314 38344
rect 12621 38335 12679 38341
rect 12621 38301 12633 38335
rect 12667 38301 12679 38335
rect 12621 38295 12679 38301
rect 10008 38236 10640 38264
rect 10008 38224 10014 38236
rect 11606 38224 11612 38276
rect 11664 38264 11670 38276
rect 12434 38264 12440 38276
rect 11664 38236 12440 38264
rect 11664 38224 11670 38236
rect 12434 38224 12440 38236
rect 12492 38264 12498 38276
rect 12636 38264 12664 38295
rect 12802 38292 12808 38344
rect 12860 38292 12866 38344
rect 12492 38236 12664 38264
rect 12492 38224 12498 38236
rect 9968 38196 9996 38224
rect 8036 38168 9996 38196
rect 12912 38196 12940 38363
rect 13633 38335 13691 38341
rect 13633 38332 13645 38335
rect 13280 38304 13645 38332
rect 13280 38273 13308 38304
rect 13633 38301 13645 38304
rect 13679 38301 13691 38335
rect 13633 38295 13691 38301
rect 15286 38292 15292 38344
rect 15344 38332 15350 38344
rect 15841 38335 15899 38341
rect 15841 38332 15853 38335
rect 15344 38304 15853 38332
rect 15344 38292 15350 38304
rect 15841 38301 15853 38304
rect 15887 38332 15899 38335
rect 15948 38332 15976 38508
rect 16485 38505 16497 38508
rect 16531 38505 16543 38539
rect 20438 38536 20444 38548
rect 16485 38499 16543 38505
rect 18064 38508 20444 38536
rect 16206 38428 16212 38480
rect 16264 38468 16270 38480
rect 18064 38468 18092 38508
rect 18138 38468 18144 38480
rect 16264 38440 17448 38468
rect 18064 38440 18144 38468
rect 16264 38428 16270 38440
rect 15887 38304 15976 38332
rect 16040 38372 16712 38400
rect 15887 38301 15899 38304
rect 15841 38295 15899 38301
rect 13265 38267 13323 38273
rect 13265 38233 13277 38267
rect 13311 38233 13323 38267
rect 13265 38227 13323 38233
rect 14642 38224 14648 38276
rect 14700 38264 14706 38276
rect 14700 38236 15240 38264
rect 14700 38224 14706 38236
rect 13998 38196 14004 38208
rect 12912 38168 14004 38196
rect 13998 38156 14004 38168
rect 14056 38156 14062 38208
rect 15102 38156 15108 38208
rect 15160 38156 15166 38208
rect 15212 38196 15240 38236
rect 16040 38196 16068 38372
rect 16390 38292 16396 38344
rect 16448 38332 16454 38344
rect 16684 38341 16712 38372
rect 17218 38360 17224 38412
rect 17276 38360 17282 38412
rect 17420 38409 17448 38440
rect 18138 38428 18144 38440
rect 18196 38428 18202 38480
rect 19812 38468 19840 38508
rect 20438 38496 20444 38508
rect 20496 38536 20502 38548
rect 20898 38536 20904 38548
rect 20496 38508 20904 38536
rect 20496 38496 20502 38508
rect 20898 38496 20904 38508
rect 20956 38496 20962 38548
rect 21082 38496 21088 38548
rect 21140 38496 21146 38548
rect 23293 38539 23351 38545
rect 23293 38505 23305 38539
rect 23339 38536 23351 38539
rect 23474 38536 23480 38548
rect 23339 38508 23480 38536
rect 23339 38505 23351 38508
rect 23293 38499 23351 38505
rect 23474 38496 23480 38508
rect 23532 38496 23538 38548
rect 23584 38508 24808 38536
rect 23584 38468 23612 38508
rect 19812 38440 20102 38468
rect 23046 38440 23612 38468
rect 23661 38471 23719 38477
rect 23661 38437 23673 38471
rect 23707 38468 23719 38471
rect 23750 38468 23756 38480
rect 23707 38440 23756 38468
rect 23707 38437 23719 38440
rect 23661 38431 23719 38437
rect 23750 38428 23756 38440
rect 23808 38428 23814 38480
rect 17405 38403 17463 38409
rect 17405 38369 17417 38403
rect 17451 38369 17463 38403
rect 17405 38363 17463 38369
rect 21542 38360 21548 38412
rect 21600 38360 21606 38412
rect 24780 38400 24808 38508
rect 25130 38496 25136 38548
rect 25188 38496 25194 38548
rect 26050 38496 26056 38548
rect 26108 38536 26114 38548
rect 27522 38536 27528 38548
rect 26108 38508 27528 38536
rect 26108 38496 26114 38508
rect 27522 38496 27528 38508
rect 27580 38496 27586 38548
rect 27614 38496 27620 38548
rect 27672 38536 27678 38548
rect 34422 38536 34428 38548
rect 27672 38508 34428 38536
rect 27672 38496 27678 38508
rect 34422 38496 34428 38508
rect 34480 38496 34486 38548
rect 34514 38496 34520 38548
rect 34572 38536 34578 38548
rect 34572 38508 34836 38536
rect 34572 38496 34578 38508
rect 29822 38428 29828 38480
rect 29880 38468 29886 38480
rect 29917 38471 29975 38477
rect 29917 38468 29929 38471
rect 29880 38440 29929 38468
rect 29880 38428 29886 38440
rect 29917 38437 29929 38440
rect 29963 38437 29975 38471
rect 30558 38468 30564 38480
rect 29917 38431 29975 38437
rect 30392 38440 30564 38468
rect 25406 38400 25412 38412
rect 24780 38386 25412 38400
rect 24794 38372 25412 38386
rect 25406 38360 25412 38372
rect 25464 38360 25470 38412
rect 26789 38403 26847 38409
rect 26789 38369 26801 38403
rect 26835 38400 26847 38403
rect 27249 38403 27307 38409
rect 27249 38400 27261 38403
rect 26835 38372 27261 38400
rect 26835 38369 26847 38372
rect 26789 38363 26847 38369
rect 27249 38369 27261 38372
rect 27295 38369 27307 38403
rect 27249 38363 27307 38369
rect 29273 38403 29331 38409
rect 29273 38369 29285 38403
rect 29319 38400 29331 38403
rect 30392 38400 30420 38440
rect 30558 38428 30564 38440
rect 30616 38428 30622 38480
rect 30742 38428 30748 38480
rect 30800 38468 30806 38480
rect 33962 38468 33968 38480
rect 30800 38440 33968 38468
rect 30800 38428 30806 38440
rect 33962 38428 33968 38440
rect 34020 38428 34026 38480
rect 34808 38468 34836 38508
rect 35434 38496 35440 38548
rect 35492 38496 35498 38548
rect 35618 38496 35624 38548
rect 35676 38536 35682 38548
rect 35805 38539 35863 38545
rect 35805 38536 35817 38539
rect 35676 38508 35817 38536
rect 35676 38496 35682 38508
rect 35805 38505 35817 38508
rect 35851 38505 35863 38539
rect 35805 38499 35863 38505
rect 38470 38496 38476 38548
rect 38528 38496 38534 38548
rect 40862 38536 40868 38548
rect 39316 38508 40868 38536
rect 35897 38471 35955 38477
rect 35897 38468 35909 38471
rect 34808 38440 35909 38468
rect 35897 38437 35909 38440
rect 35943 38437 35955 38471
rect 35897 38431 35955 38437
rect 36998 38428 37004 38480
rect 37056 38428 37062 38480
rect 29319 38372 30420 38400
rect 29319 38369 29331 38372
rect 29273 38363 29331 38369
rect 30466 38360 30472 38412
rect 30524 38360 30530 38412
rect 31021 38403 31079 38409
rect 31021 38369 31033 38403
rect 31067 38400 31079 38403
rect 31386 38400 31392 38412
rect 31067 38372 31392 38400
rect 31067 38369 31079 38372
rect 31021 38363 31079 38369
rect 16577 38335 16635 38341
rect 16577 38332 16589 38335
rect 16448 38304 16589 38332
rect 16448 38292 16454 38304
rect 16577 38301 16589 38304
rect 16623 38301 16635 38335
rect 16577 38295 16635 38301
rect 16669 38335 16727 38341
rect 16669 38301 16681 38335
rect 16715 38301 16727 38335
rect 16669 38295 16727 38301
rect 16592 38264 16620 38295
rect 17678 38292 17684 38344
rect 17736 38292 17742 38344
rect 19334 38292 19340 38344
rect 19392 38292 19398 38344
rect 19613 38335 19671 38341
rect 19613 38301 19625 38335
rect 19659 38332 19671 38335
rect 20254 38332 20260 38344
rect 19659 38304 20260 38332
rect 19659 38301 19671 38304
rect 19613 38295 19671 38301
rect 20254 38292 20260 38304
rect 20312 38292 20318 38344
rect 21821 38335 21879 38341
rect 21821 38301 21833 38335
rect 21867 38332 21879 38335
rect 22830 38332 22836 38344
rect 21867 38304 22836 38332
rect 21867 38301 21879 38304
rect 21821 38295 21879 38301
rect 22830 38292 22836 38304
rect 22888 38292 22894 38344
rect 23385 38335 23443 38341
rect 23385 38332 23397 38335
rect 23308 38304 23397 38332
rect 23308 38264 23336 38304
rect 23385 38301 23397 38304
rect 23431 38301 23443 38335
rect 23658 38332 23664 38344
rect 23385 38295 23443 38301
rect 23492 38304 23664 38332
rect 23492 38264 23520 38304
rect 23658 38292 23664 38304
rect 23716 38332 23722 38344
rect 26142 38332 26148 38344
rect 23716 38304 26148 38332
rect 23716 38292 23722 38304
rect 26142 38292 26148 38304
rect 26200 38292 26206 38344
rect 26878 38292 26884 38344
rect 26936 38292 26942 38344
rect 26973 38335 27031 38341
rect 26973 38301 26985 38335
rect 27019 38301 27031 38335
rect 26973 38295 27031 38301
rect 16592 38236 16712 38264
rect 23308 38236 23520 38264
rect 15212 38168 16068 38196
rect 16114 38156 16120 38208
rect 16172 38156 16178 38208
rect 16684 38196 16712 38236
rect 23492 38208 23520 38236
rect 26234 38224 26240 38276
rect 26292 38264 26298 38276
rect 26292 38236 26740 38264
rect 26292 38224 26298 38236
rect 19058 38196 19064 38208
rect 16684 38168 19064 38196
rect 19058 38156 19064 38168
rect 19116 38156 19122 38208
rect 19153 38199 19211 38205
rect 19153 38165 19165 38199
rect 19199 38196 19211 38199
rect 19242 38196 19248 38208
rect 19199 38168 19248 38196
rect 19199 38165 19211 38168
rect 19153 38159 19211 38165
rect 19242 38156 19248 38168
rect 19300 38156 19306 38208
rect 23474 38156 23480 38208
rect 23532 38156 23538 38208
rect 25682 38156 25688 38208
rect 25740 38196 25746 38208
rect 26421 38199 26479 38205
rect 26421 38196 26433 38199
rect 25740 38168 26433 38196
rect 25740 38156 25746 38168
rect 26421 38165 26433 38168
rect 26467 38165 26479 38199
rect 26712 38196 26740 38236
rect 26786 38224 26792 38276
rect 26844 38264 26850 38276
rect 26988 38264 27016 38295
rect 27798 38292 27804 38344
rect 27856 38292 27862 38344
rect 29178 38292 29184 38344
rect 29236 38332 29242 38344
rect 29365 38335 29423 38341
rect 29365 38332 29377 38335
rect 29236 38304 29377 38332
rect 29236 38292 29242 38304
rect 29365 38301 29377 38304
rect 29411 38301 29423 38335
rect 29365 38295 29423 38301
rect 29457 38335 29515 38341
rect 29457 38301 29469 38335
rect 29503 38301 29515 38335
rect 29457 38295 29515 38301
rect 26844 38236 27016 38264
rect 26844 38224 26850 38236
rect 28166 38224 28172 38276
rect 28224 38264 28230 38276
rect 28905 38267 28963 38273
rect 28905 38264 28917 38267
rect 28224 38236 28917 38264
rect 28224 38224 28230 38236
rect 28905 38233 28917 38236
rect 28951 38233 28963 38267
rect 28905 38227 28963 38233
rect 28626 38196 28632 38208
rect 26712 38168 28632 38196
rect 26421 38159 26479 38165
rect 28626 38156 28632 38168
rect 28684 38196 28690 38208
rect 29472 38196 29500 38295
rect 30006 38292 30012 38344
rect 30064 38332 30070 38344
rect 31036 38332 31064 38363
rect 31386 38360 31392 38372
rect 31444 38400 31450 38412
rect 31573 38403 31631 38409
rect 31573 38400 31585 38403
rect 31444 38372 31585 38400
rect 31444 38360 31450 38372
rect 31573 38369 31585 38372
rect 31619 38369 31631 38403
rect 31573 38363 31631 38369
rect 33134 38360 33140 38412
rect 33192 38400 33198 38412
rect 33229 38403 33287 38409
rect 33229 38400 33241 38403
rect 33192 38372 33241 38400
rect 33192 38360 33198 38372
rect 33229 38369 33241 38372
rect 33275 38369 33287 38403
rect 36449 38403 36507 38409
rect 36449 38400 36461 38403
rect 33229 38363 33287 38369
rect 34992 38372 36461 38400
rect 30064 38304 31064 38332
rect 30064 38292 30070 38304
rect 31110 38292 31116 38344
rect 31168 38292 31174 38344
rect 31297 38335 31355 38341
rect 31297 38301 31309 38335
rect 31343 38332 31355 38335
rect 31478 38332 31484 38344
rect 31343 38304 31484 38332
rect 31343 38301 31355 38304
rect 31297 38295 31355 38301
rect 31478 38292 31484 38304
rect 31536 38292 31542 38344
rect 33505 38335 33563 38341
rect 33505 38301 33517 38335
rect 33551 38332 33563 38335
rect 34238 38332 34244 38344
rect 33551 38304 34244 38332
rect 33551 38301 33563 38304
rect 33505 38295 33563 38301
rect 34238 38292 34244 38304
rect 34296 38292 34302 38344
rect 34698 38292 34704 38344
rect 34756 38332 34762 38344
rect 34992 38341 35020 38372
rect 36449 38369 36461 38372
rect 36495 38369 36507 38403
rect 36449 38363 36507 38369
rect 36722 38360 36728 38412
rect 36780 38360 36786 38412
rect 39316 38409 39344 38508
rect 40862 38496 40868 38508
rect 40920 38496 40926 38548
rect 41414 38496 41420 38548
rect 41472 38536 41478 38548
rect 41877 38539 41935 38545
rect 41877 38536 41889 38539
rect 41472 38508 41889 38536
rect 41472 38496 41478 38508
rect 41877 38505 41889 38508
rect 41923 38505 41935 38539
rect 41877 38499 41935 38505
rect 42337 38539 42395 38545
rect 42337 38505 42349 38539
rect 42383 38536 42395 38539
rect 42610 38536 42616 38548
rect 42383 38508 42616 38536
rect 42383 38505 42395 38508
rect 42337 38499 42395 38505
rect 42610 38496 42616 38508
rect 42668 38496 42674 38548
rect 42702 38496 42708 38548
rect 42760 38536 42766 38548
rect 42760 38508 44680 38536
rect 42760 38496 42766 38508
rect 39577 38471 39635 38477
rect 39577 38437 39589 38471
rect 39623 38468 39635 38471
rect 39850 38468 39856 38480
rect 39623 38440 39856 38468
rect 39623 38437 39635 38440
rect 39577 38431 39635 38437
rect 39850 38428 39856 38440
rect 39908 38428 39914 38480
rect 40034 38428 40040 38480
rect 40092 38428 40098 38480
rect 44542 38428 44548 38480
rect 44600 38428 44606 38480
rect 44652 38468 44680 38508
rect 45186 38496 45192 38548
rect 45244 38536 45250 38548
rect 45373 38539 45431 38545
rect 45373 38536 45385 38539
rect 45244 38508 45385 38536
rect 45244 38496 45250 38508
rect 45373 38505 45385 38508
rect 45419 38505 45431 38539
rect 45373 38499 45431 38505
rect 46109 38539 46167 38545
rect 46109 38505 46121 38539
rect 46155 38536 46167 38539
rect 46198 38536 46204 38548
rect 46155 38508 46204 38536
rect 46155 38505 46167 38508
rect 46109 38499 46167 38505
rect 46198 38496 46204 38508
rect 46256 38496 46262 38548
rect 46477 38539 46535 38545
rect 46477 38505 46489 38539
rect 46523 38536 46535 38539
rect 47762 38536 47768 38548
rect 46523 38508 47768 38536
rect 46523 38505 46535 38508
rect 46477 38499 46535 38505
rect 47762 38496 47768 38508
rect 47820 38496 47826 38548
rect 47872 38508 50292 38536
rect 47872 38468 47900 38508
rect 44652 38440 47900 38468
rect 48958 38428 48964 38480
rect 49016 38428 49022 38480
rect 49694 38428 49700 38480
rect 49752 38428 49758 38480
rect 50264 38468 50292 38508
rect 50338 38496 50344 38548
rect 50396 38536 50402 38548
rect 50433 38539 50491 38545
rect 50433 38536 50445 38539
rect 50396 38508 50445 38536
rect 50396 38496 50402 38508
rect 50433 38505 50445 38508
rect 50479 38505 50491 38539
rect 50433 38499 50491 38505
rect 50982 38496 50988 38548
rect 51040 38496 51046 38548
rect 63770 38536 63776 38548
rect 53576 38508 63776 38536
rect 53576 38468 53604 38508
rect 63770 38496 63776 38508
rect 63828 38496 63834 38548
rect 50264 38440 53604 38468
rect 53834 38428 53840 38480
rect 53892 38428 53898 38480
rect 55493 38471 55551 38477
rect 55493 38437 55505 38471
rect 55539 38468 55551 38471
rect 55766 38468 55772 38480
rect 55539 38440 55772 38468
rect 55539 38437 55551 38440
rect 55493 38431 55551 38437
rect 55766 38428 55772 38440
rect 55824 38428 55830 38480
rect 55950 38428 55956 38480
rect 56008 38428 56014 38480
rect 58342 38428 58348 38480
rect 58400 38468 58406 38480
rect 58400 38440 58558 38468
rect 58400 38428 58406 38440
rect 60734 38428 60740 38480
rect 60792 38468 60798 38480
rect 62482 38468 62488 38480
rect 60792 38440 62488 38468
rect 60792 38428 60798 38440
rect 62482 38428 62488 38440
rect 62540 38428 62546 38480
rect 39301 38403 39359 38409
rect 34977 38335 35035 38341
rect 34977 38332 34989 38335
rect 34756 38304 34989 38332
rect 34756 38292 34762 38304
rect 34977 38301 34989 38304
rect 35023 38301 35035 38335
rect 34977 38295 35035 38301
rect 35158 38292 35164 38344
rect 35216 38292 35222 38344
rect 35250 38292 35256 38344
rect 35308 38332 35314 38344
rect 35345 38335 35403 38341
rect 35345 38332 35357 38335
rect 35308 38304 35357 38332
rect 35308 38292 35314 38304
rect 35345 38301 35357 38304
rect 35391 38301 35403 38335
rect 38120 38332 38148 38386
rect 39301 38369 39313 38403
rect 39347 38369 39359 38403
rect 39301 38363 39359 38369
rect 40862 38360 40868 38412
rect 40920 38400 40926 38412
rect 41322 38400 41328 38412
rect 40920 38372 41328 38400
rect 40920 38360 40926 38372
rect 41322 38360 41328 38372
rect 41380 38360 41386 38412
rect 42245 38403 42303 38409
rect 42245 38369 42257 38403
rect 42291 38400 42303 38403
rect 42705 38403 42763 38409
rect 42705 38400 42717 38403
rect 42291 38372 42717 38400
rect 42291 38369 42303 38372
rect 42245 38363 42303 38369
rect 42705 38369 42717 38372
rect 42751 38369 42763 38403
rect 42705 38363 42763 38369
rect 43254 38360 43260 38412
rect 43312 38360 43318 38412
rect 45278 38360 45284 38412
rect 45336 38360 45342 38412
rect 47302 38400 47308 38412
rect 46676 38372 47308 38400
rect 38746 38332 38752 38344
rect 38120 38304 38752 38332
rect 35345 38295 35403 38301
rect 38746 38292 38752 38304
rect 38804 38332 38810 38344
rect 39942 38332 39948 38344
rect 38804 38304 39948 38332
rect 38804 38292 38810 38304
rect 39942 38292 39948 38304
rect 40000 38292 40006 38344
rect 40770 38292 40776 38344
rect 40828 38332 40834 38344
rect 41598 38332 41604 38344
rect 40828 38304 41604 38332
rect 40828 38292 40834 38304
rect 41598 38292 41604 38304
rect 41656 38292 41662 38344
rect 42518 38292 42524 38344
rect 42576 38292 42582 38344
rect 44450 38292 44456 38344
rect 44508 38332 44514 38344
rect 45005 38335 45063 38341
rect 45005 38332 45017 38335
rect 44508 38304 45017 38332
rect 44508 38292 44514 38304
rect 45005 38301 45017 38304
rect 45051 38301 45063 38335
rect 45005 38295 45063 38301
rect 45925 38335 45983 38341
rect 45925 38301 45937 38335
rect 45971 38301 45983 38335
rect 45925 38295 45983 38301
rect 29546 38224 29552 38276
rect 29604 38264 29610 38276
rect 41506 38264 41512 38276
rect 29604 38236 33364 38264
rect 29604 38224 29610 38236
rect 28684 38168 29500 38196
rect 28684 38156 28690 38168
rect 30650 38156 30656 38208
rect 30708 38156 30714 38208
rect 32214 38156 32220 38208
rect 32272 38156 32278 38208
rect 33336 38196 33364 38236
rect 34624 38236 36584 38264
rect 34624 38196 34652 38236
rect 33336 38168 34652 38196
rect 36556 38196 36584 38236
rect 38028 38236 38608 38264
rect 38028 38196 38056 38236
rect 36556 38168 38056 38196
rect 38580 38196 38608 38236
rect 40604 38236 41512 38264
rect 40604 38196 40632 38236
rect 41506 38224 41512 38236
rect 41564 38224 41570 38276
rect 43990 38264 43996 38276
rect 43456 38236 43996 38264
rect 38580 38168 40632 38196
rect 40770 38156 40776 38208
rect 40828 38196 40834 38208
rect 41049 38199 41107 38205
rect 41049 38196 41061 38199
rect 40828 38168 41061 38196
rect 40828 38156 40834 38168
rect 41049 38165 41061 38168
rect 41095 38165 41107 38199
rect 41049 38159 41107 38165
rect 41322 38156 41328 38208
rect 41380 38196 41386 38208
rect 43456 38196 43484 38236
rect 43990 38224 43996 38236
rect 44048 38224 44054 38276
rect 41380 38168 43484 38196
rect 43533 38199 43591 38205
rect 41380 38156 41386 38168
rect 43533 38165 43545 38199
rect 43579 38196 43591 38199
rect 43806 38196 43812 38208
rect 43579 38168 43812 38196
rect 43579 38165 43591 38168
rect 43533 38159 43591 38165
rect 43806 38156 43812 38168
rect 43864 38156 43870 38208
rect 44818 38156 44824 38208
rect 44876 38196 44882 38208
rect 45940 38196 45968 38295
rect 46566 38292 46572 38344
rect 46624 38292 46630 38344
rect 46676 38341 46704 38372
rect 47302 38360 47308 38372
rect 47360 38400 47366 38412
rect 47670 38400 47676 38412
rect 47360 38372 47676 38400
rect 47360 38360 47366 38372
rect 47670 38360 47676 38372
rect 47728 38360 47734 38412
rect 48222 38360 48228 38412
rect 48280 38400 48286 38412
rect 48685 38403 48743 38409
rect 48685 38400 48697 38403
rect 48280 38372 48697 38400
rect 48280 38360 48286 38372
rect 48685 38369 48697 38372
rect 48731 38369 48743 38403
rect 48685 38363 48743 38369
rect 50798 38360 50804 38412
rect 50856 38400 50862 38412
rect 64966 38400 64972 38412
rect 50856 38372 51212 38400
rect 50856 38360 50862 38372
rect 46661 38335 46719 38341
rect 46661 38301 46673 38335
rect 46707 38301 46719 38335
rect 46661 38295 46719 38301
rect 46750 38292 46756 38344
rect 46808 38332 46814 38344
rect 47029 38335 47087 38341
rect 47029 38332 47041 38335
rect 46808 38304 47041 38332
rect 46808 38292 46814 38304
rect 47029 38301 47041 38304
rect 47075 38301 47087 38335
rect 47029 38295 47087 38301
rect 50890 38292 50896 38344
rect 50948 38332 50954 38344
rect 51184 38341 51212 38372
rect 59096 38372 64972 38400
rect 51077 38335 51135 38341
rect 51077 38332 51089 38335
rect 50948 38304 51089 38332
rect 50948 38292 50954 38304
rect 51077 38301 51089 38304
rect 51123 38301 51135 38335
rect 51077 38295 51135 38301
rect 51169 38335 51227 38341
rect 51169 38301 51181 38335
rect 51215 38301 51227 38335
rect 51169 38295 51227 38301
rect 51718 38292 51724 38344
rect 51776 38332 51782 38344
rect 52733 38335 52791 38341
rect 52733 38332 52745 38335
rect 51776 38304 52745 38332
rect 51776 38292 51782 38304
rect 52733 38301 52745 38304
rect 52779 38301 52791 38335
rect 52733 38295 52791 38301
rect 53101 38335 53159 38341
rect 53101 38301 53113 38335
rect 53147 38332 53159 38335
rect 54110 38332 54116 38344
rect 53147 38304 54116 38332
rect 53147 38301 53159 38304
rect 53101 38295 53159 38301
rect 49970 38224 49976 38276
rect 50028 38264 50034 38276
rect 53116 38264 53144 38295
rect 54110 38292 54116 38304
rect 54168 38292 54174 38344
rect 54386 38292 54392 38344
rect 54444 38332 54450 38344
rect 54849 38335 54907 38341
rect 54849 38332 54861 38335
rect 54444 38304 54861 38332
rect 54444 38292 54450 38304
rect 54849 38301 54861 38304
rect 54895 38301 54907 38335
rect 54849 38295 54907 38301
rect 55125 38335 55183 38341
rect 55125 38301 55137 38335
rect 55171 38301 55183 38335
rect 55125 38295 55183 38301
rect 50028 38236 53144 38264
rect 55140 38264 55168 38295
rect 55214 38292 55220 38344
rect 55272 38292 55278 38344
rect 57790 38332 57796 38344
rect 55324 38304 57796 38332
rect 55324 38264 55352 38304
rect 57790 38292 57796 38304
rect 57848 38292 57854 38344
rect 58069 38335 58127 38341
rect 58069 38301 58081 38335
rect 58115 38332 58127 38335
rect 58158 38332 58164 38344
rect 58115 38304 58164 38332
rect 58115 38301 58127 38304
rect 58069 38295 58127 38301
rect 58158 38292 58164 38304
rect 58216 38292 58222 38344
rect 58434 38292 58440 38344
rect 58492 38332 58498 38344
rect 59096 38332 59124 38372
rect 64966 38360 64972 38372
rect 65024 38360 65030 38412
rect 58492 38304 59124 38332
rect 58492 38292 58498 38304
rect 59262 38292 59268 38344
rect 59320 38332 59326 38344
rect 59817 38335 59875 38341
rect 59817 38332 59829 38335
rect 59320 38304 59829 38332
rect 59320 38292 59326 38304
rect 59817 38301 59829 38304
rect 59863 38301 59875 38335
rect 59817 38295 59875 38301
rect 55140 38236 55352 38264
rect 50028 38224 50034 38236
rect 56778 38224 56784 38276
rect 56836 38264 56842 38276
rect 56836 38236 57836 38264
rect 56836 38224 56842 38236
rect 44876 38168 45968 38196
rect 44876 38156 44882 38168
rect 47486 38156 47492 38208
rect 47544 38196 47550 38208
rect 47673 38199 47731 38205
rect 47673 38196 47685 38199
rect 47544 38168 47685 38196
rect 47544 38156 47550 38168
rect 47673 38165 47685 38168
rect 47719 38165 47731 38199
rect 47673 38159 47731 38165
rect 50614 38156 50620 38208
rect 50672 38156 50678 38208
rect 51626 38156 51632 38208
rect 51684 38196 51690 38208
rect 52181 38199 52239 38205
rect 52181 38196 52193 38199
rect 51684 38168 52193 38196
rect 51684 38156 51690 38168
rect 52181 38165 52193 38168
rect 52227 38165 52239 38199
rect 52181 38159 52239 38165
rect 56965 38199 57023 38205
rect 56965 38165 56977 38199
rect 57011 38196 57023 38199
rect 57146 38196 57152 38208
rect 57011 38168 57152 38196
rect 57011 38165 57023 38168
rect 56965 38159 57023 38165
rect 57146 38156 57152 38168
rect 57204 38196 57210 38208
rect 57698 38196 57704 38208
rect 57204 38168 57704 38196
rect 57204 38156 57210 38168
rect 57698 38156 57704 38168
rect 57756 38156 57762 38208
rect 57808 38196 57836 38236
rect 63310 38196 63316 38208
rect 57808 38168 63316 38196
rect 63310 38156 63316 38168
rect 63368 38156 63374 38208
rect 552 38106 66424 38128
rect 552 38054 1998 38106
rect 2050 38054 2062 38106
rect 2114 38054 2126 38106
rect 2178 38054 2190 38106
rect 2242 38054 2254 38106
rect 2306 38054 50998 38106
rect 51050 38054 51062 38106
rect 51114 38054 51126 38106
rect 51178 38054 51190 38106
rect 51242 38054 51254 38106
rect 51306 38054 66424 38106
rect 552 38032 66424 38054
rect 7374 37952 7380 38004
rect 7432 37992 7438 38004
rect 9585 37995 9643 38001
rect 9585 37992 9597 37995
rect 7432 37964 9597 37992
rect 7432 37952 7438 37964
rect 9585 37961 9597 37964
rect 9631 37961 9643 37995
rect 9585 37955 9643 37961
rect 9858 37952 9864 38004
rect 9916 37992 9922 38004
rect 10413 37995 10471 38001
rect 10413 37992 10425 37995
rect 9916 37964 10425 37992
rect 9916 37952 9922 37964
rect 10413 37961 10425 37964
rect 10459 37961 10471 37995
rect 10413 37955 10471 37961
rect 14277 37995 14335 38001
rect 14277 37961 14289 37995
rect 14323 37992 14335 37995
rect 15378 37992 15384 38004
rect 14323 37964 15384 37992
rect 14323 37961 14335 37964
rect 14277 37955 14335 37961
rect 15378 37952 15384 37964
rect 15436 37952 15442 38004
rect 15767 37995 15825 38001
rect 15767 37961 15779 37995
rect 15813 37992 15825 37995
rect 16114 37992 16120 38004
rect 15813 37964 16120 37992
rect 15813 37961 15825 37964
rect 15767 37955 15825 37961
rect 16114 37952 16120 37964
rect 16172 37952 16178 38004
rect 17218 37952 17224 38004
rect 17276 37992 17282 38004
rect 19334 37992 19340 38004
rect 17276 37964 19340 37992
rect 17276 37952 17282 37964
rect 19334 37952 19340 37964
rect 19392 37992 19398 38004
rect 24660 37995 24718 38001
rect 19392 37964 24440 37992
rect 19392 37952 19398 37964
rect 7926 37884 7932 37936
rect 7984 37924 7990 37936
rect 12434 37924 12440 37936
rect 7984 37896 12440 37924
rect 7984 37884 7990 37896
rect 6457 37859 6515 37865
rect 6457 37825 6469 37859
rect 6503 37856 6515 37859
rect 7098 37856 7104 37868
rect 6503 37828 7104 37856
rect 6503 37825 6515 37828
rect 6457 37819 6515 37825
rect 7098 37816 7104 37828
rect 7156 37816 7162 37868
rect 9416 37865 9444 37896
rect 12434 37884 12440 37896
rect 12492 37924 12498 37936
rect 14642 37924 14648 37936
rect 12492 37896 14648 37924
rect 12492 37884 12498 37896
rect 14642 37884 14648 37896
rect 14700 37884 14706 37936
rect 18046 37884 18052 37936
rect 18104 37924 18110 37936
rect 18693 37927 18751 37933
rect 18693 37924 18705 37927
rect 18104 37896 18705 37924
rect 18104 37884 18110 37896
rect 18693 37893 18705 37896
rect 18739 37893 18751 37927
rect 18693 37887 18751 37893
rect 22830 37884 22836 37936
rect 22888 37924 22894 37936
rect 22925 37927 22983 37933
rect 22925 37924 22937 37927
rect 22888 37896 22937 37924
rect 22888 37884 22894 37896
rect 22925 37893 22937 37896
rect 22971 37893 22983 37927
rect 22925 37887 22983 37893
rect 23290 37884 23296 37936
rect 23348 37924 23354 37936
rect 23348 37896 23520 37924
rect 23348 37884 23354 37896
rect 8205 37859 8263 37865
rect 8205 37825 8217 37859
rect 8251 37825 8263 37859
rect 8205 37819 8263 37825
rect 9401 37859 9459 37865
rect 9401 37825 9413 37859
rect 9447 37825 9459 37859
rect 9401 37819 9459 37825
rect 10229 37859 10287 37865
rect 10229 37825 10241 37859
rect 10275 37856 10287 37859
rect 10965 37859 11023 37865
rect 10965 37856 10977 37859
rect 10275 37828 10977 37856
rect 10275 37825 10287 37828
rect 10229 37819 10287 37825
rect 10965 37825 10977 37828
rect 11011 37856 11023 37859
rect 12250 37856 12256 37868
rect 11011 37828 12256 37856
rect 11011 37825 11023 37828
rect 10965 37819 11023 37825
rect 8220 37788 8248 37819
rect 12250 37816 12256 37828
rect 12308 37816 12314 37868
rect 12802 37816 12808 37868
rect 12860 37856 12866 37868
rect 15102 37856 15108 37868
rect 12860 37828 15108 37856
rect 12860 37816 12866 37828
rect 15102 37816 15108 37828
rect 15160 37816 15166 37868
rect 15194 37816 15200 37868
rect 15252 37856 15258 37868
rect 16025 37859 16083 37865
rect 16025 37856 16037 37859
rect 15252 37828 16037 37856
rect 15252 37816 15258 37828
rect 16025 37825 16037 37828
rect 16071 37825 16083 37859
rect 16025 37819 16083 37825
rect 19245 37859 19303 37865
rect 19245 37825 19257 37859
rect 19291 37856 19303 37859
rect 20533 37859 20591 37865
rect 19291 37828 20484 37856
rect 19291 37825 19303 37828
rect 19245 37819 19303 37825
rect 9125 37791 9183 37797
rect 9125 37788 9137 37791
rect 8220 37760 9137 37788
rect 9125 37757 9137 37760
rect 9171 37788 9183 37791
rect 11514 37788 11520 37800
rect 9171 37760 11520 37788
rect 9171 37757 9183 37760
rect 9125 37751 9183 37757
rect 11514 37748 11520 37760
rect 11572 37748 11578 37800
rect 14274 37748 14280 37800
rect 14332 37788 14338 37800
rect 16040 37788 16068 37819
rect 16206 37788 16212 37800
rect 14332 37760 14674 37788
rect 16040 37760 16212 37788
rect 14332 37748 14338 37760
rect 16206 37748 16212 37760
rect 16264 37748 16270 37800
rect 18509 37791 18567 37797
rect 18509 37757 18521 37791
rect 18555 37788 18567 37791
rect 18690 37788 18696 37800
rect 18555 37760 18696 37788
rect 18555 37757 18567 37760
rect 18509 37751 18567 37757
rect 18690 37748 18696 37760
rect 18748 37748 18754 37800
rect 19150 37748 19156 37800
rect 19208 37748 19214 37800
rect 6733 37723 6791 37729
rect 6733 37689 6745 37723
rect 6779 37720 6791 37723
rect 7006 37720 7012 37732
rect 6779 37692 7012 37720
rect 6779 37689 6791 37692
rect 6733 37683 6791 37689
rect 7006 37680 7012 37692
rect 7064 37680 7070 37732
rect 9030 37720 9036 37732
rect 7958 37692 9036 37720
rect 9030 37680 9036 37692
rect 9088 37680 9094 37732
rect 9217 37723 9275 37729
rect 9217 37689 9229 37723
rect 9263 37720 9275 37723
rect 10873 37723 10931 37729
rect 9263 37692 10088 37720
rect 9263 37689 9275 37692
rect 9217 37683 9275 37689
rect 8754 37612 8760 37664
rect 8812 37612 8818 37664
rect 9950 37612 9956 37664
rect 10008 37612 10014 37664
rect 10060 37661 10088 37692
rect 10873 37689 10885 37723
rect 10919 37720 10931 37723
rect 12066 37720 12072 37732
rect 10919 37692 12072 37720
rect 10919 37689 10931 37692
rect 10873 37683 10931 37689
rect 12066 37680 12072 37692
rect 12124 37680 12130 37732
rect 19061 37723 19119 37729
rect 19061 37689 19073 37723
rect 19107 37720 19119 37723
rect 19242 37720 19248 37732
rect 19107 37692 19248 37720
rect 19107 37689 19119 37692
rect 19061 37683 19119 37689
rect 19242 37680 19248 37692
rect 19300 37680 19306 37732
rect 20456 37720 20484 37828
rect 20533 37825 20545 37859
rect 20579 37856 20591 37859
rect 23382 37856 23388 37868
rect 20579 37828 23388 37856
rect 20579 37825 20591 37828
rect 20533 37819 20591 37825
rect 23382 37816 23388 37828
rect 23440 37816 23446 37868
rect 23492 37865 23520 37896
rect 24412 37865 24440 37964
rect 24660 37961 24672 37995
rect 24706 37992 24718 37995
rect 25682 37992 25688 38004
rect 24706 37964 25688 37992
rect 24706 37961 24718 37964
rect 24660 37955 24718 37961
rect 25682 37952 25688 37964
rect 25740 37952 25746 38004
rect 26878 37952 26884 38004
rect 26936 37992 26942 38004
rect 28077 37995 28135 38001
rect 28077 37992 28089 37995
rect 26936 37964 28089 37992
rect 26936 37952 26942 37964
rect 28077 37961 28089 37964
rect 28123 37961 28135 37995
rect 28077 37955 28135 37961
rect 28184 37964 44128 37992
rect 25976 37896 26372 37924
rect 23477 37859 23535 37865
rect 23477 37825 23489 37859
rect 23523 37825 23535 37859
rect 23477 37819 23535 37825
rect 24397 37859 24455 37865
rect 24397 37825 24409 37859
rect 24443 37825 24455 37859
rect 24397 37819 24455 37825
rect 23014 37748 23020 37800
rect 23072 37788 23078 37800
rect 23293 37791 23351 37797
rect 23293 37788 23305 37791
rect 23072 37760 23305 37788
rect 23072 37748 23078 37760
rect 23293 37757 23305 37760
rect 23339 37757 23351 37791
rect 23293 37751 23351 37757
rect 20714 37720 20720 37732
rect 20456 37692 20720 37720
rect 20714 37680 20720 37692
rect 20772 37680 20778 37732
rect 20806 37680 20812 37732
rect 20864 37680 20870 37732
rect 20898 37680 20904 37732
rect 20956 37720 20962 37732
rect 20956 37692 21298 37720
rect 22204 37692 23980 37720
rect 20956 37680 20962 37692
rect 10045 37655 10103 37661
rect 10045 37621 10057 37655
rect 10091 37652 10103 37655
rect 10502 37652 10508 37664
rect 10091 37624 10508 37652
rect 10091 37621 10103 37624
rect 10045 37615 10103 37621
rect 10502 37612 10508 37624
rect 10560 37652 10566 37664
rect 10781 37655 10839 37661
rect 10781 37652 10793 37655
rect 10560 37624 10793 37652
rect 10560 37612 10566 37624
rect 10781 37621 10793 37624
rect 10827 37621 10839 37655
rect 10781 37615 10839 37621
rect 15010 37612 15016 37664
rect 15068 37652 15074 37664
rect 22204 37652 22232 37692
rect 15068 37624 22232 37652
rect 15068 37612 15074 37624
rect 22278 37612 22284 37664
rect 22336 37612 22342 37664
rect 23385 37655 23443 37661
rect 23385 37621 23397 37655
rect 23431 37652 23443 37655
rect 23842 37652 23848 37664
rect 23431 37624 23848 37652
rect 23431 37621 23443 37624
rect 23385 37615 23443 37621
rect 23842 37612 23848 37624
rect 23900 37612 23906 37664
rect 23952 37652 23980 37692
rect 25406 37680 25412 37732
rect 25464 37680 25470 37732
rect 25976 37652 26004 37896
rect 26142 37816 26148 37868
rect 26200 37856 26206 37868
rect 26237 37859 26295 37865
rect 26237 37856 26249 37859
rect 26200 37828 26249 37856
rect 26200 37816 26206 37828
rect 26237 37825 26249 37828
rect 26283 37825 26295 37859
rect 26344 37856 26372 37896
rect 27614 37884 27620 37936
rect 27672 37924 27678 37936
rect 27982 37924 27988 37936
rect 27672 37896 27988 37924
rect 27672 37884 27678 37896
rect 27982 37884 27988 37896
rect 28040 37884 28046 37936
rect 28184 37856 28212 37964
rect 30650 37924 30656 37936
rect 29932 37896 30656 37924
rect 26344 37828 28212 37856
rect 26237 37819 26295 37825
rect 28626 37816 28632 37868
rect 28684 37816 28690 37868
rect 29932 37865 29960 37896
rect 30650 37884 30656 37896
rect 30708 37884 30714 37936
rect 31956 37896 32812 37924
rect 29917 37859 29975 37865
rect 29917 37825 29929 37859
rect 29963 37825 29975 37859
rect 29917 37819 29975 37825
rect 30101 37859 30159 37865
rect 30101 37825 30113 37859
rect 30147 37856 30159 37859
rect 30282 37856 30288 37868
rect 30147 37828 30288 37856
rect 30147 37825 30159 37828
rect 30101 37819 30159 37825
rect 30282 37816 30288 37828
rect 30340 37816 30346 37868
rect 31956 37856 31984 37896
rect 30576 37828 31984 37856
rect 27614 37748 27620 37800
rect 27672 37748 27678 37800
rect 27890 37748 27896 37800
rect 27948 37788 27954 37800
rect 30576 37788 30604 37828
rect 32030 37816 32036 37868
rect 32088 37816 32094 37868
rect 27948 37760 30604 37788
rect 27948 37748 27954 37760
rect 30650 37748 30656 37800
rect 30708 37748 30714 37800
rect 32677 37791 32735 37797
rect 32677 37757 32689 37791
rect 32723 37757 32735 37791
rect 32677 37751 32735 37757
rect 26510 37680 26516 37732
rect 26568 37680 26574 37732
rect 28445 37723 28503 37729
rect 28445 37720 28457 37723
rect 28000 37692 28457 37720
rect 23952 37624 26004 37652
rect 26145 37655 26203 37661
rect 26145 37621 26157 37655
rect 26191 37652 26203 37655
rect 27798 37652 27804 37664
rect 26191 37624 27804 37652
rect 26191 37621 26203 37624
rect 26145 37615 26203 37621
rect 27798 37612 27804 37624
rect 27856 37612 27862 37664
rect 28000 37661 28028 37692
rect 28445 37689 28457 37692
rect 28491 37720 28503 37723
rect 29178 37720 29184 37732
rect 28491 37692 29184 37720
rect 28491 37689 28503 37692
rect 28445 37683 28503 37689
rect 29178 37680 29184 37692
rect 29236 37680 29242 37732
rect 29825 37723 29883 37729
rect 29825 37689 29837 37723
rect 29871 37720 29883 37723
rect 29871 37692 30512 37720
rect 29871 37689 29883 37692
rect 29825 37683 29883 37689
rect 27985 37655 28043 37661
rect 27985 37621 27997 37655
rect 28031 37621 28043 37655
rect 27985 37615 28043 37621
rect 28534 37612 28540 37664
rect 28592 37612 28598 37664
rect 29457 37655 29515 37661
rect 29457 37621 29469 37655
rect 29503 37652 29515 37655
rect 29638 37652 29644 37664
rect 29503 37624 29644 37652
rect 29503 37621 29515 37624
rect 29457 37615 29515 37621
rect 29638 37612 29644 37624
rect 29696 37612 29702 37664
rect 30006 37612 30012 37664
rect 30064 37652 30070 37664
rect 30285 37655 30343 37661
rect 30285 37652 30297 37655
rect 30064 37624 30297 37652
rect 30064 37612 30070 37624
rect 30285 37621 30297 37624
rect 30331 37621 30343 37655
rect 30484 37652 30512 37692
rect 31662 37680 31668 37732
rect 31720 37720 31726 37732
rect 31757 37723 31815 37729
rect 31757 37720 31769 37723
rect 31720 37692 31769 37720
rect 31720 37680 31726 37692
rect 31757 37689 31769 37692
rect 31803 37689 31815 37723
rect 31757 37683 31815 37689
rect 31846 37680 31852 37732
rect 31904 37720 31910 37732
rect 32692 37720 32720 37751
rect 31904 37692 32720 37720
rect 32784 37720 32812 37896
rect 34238 37884 34244 37936
rect 34296 37884 34302 37936
rect 34330 37884 34336 37936
rect 34388 37924 34394 37936
rect 34388 37896 37320 37924
rect 34388 37884 34394 37896
rect 34885 37859 34943 37865
rect 34885 37825 34897 37859
rect 34931 37856 34943 37859
rect 35158 37856 35164 37868
rect 34931 37828 35164 37856
rect 34931 37825 34943 37828
rect 34885 37819 34943 37825
rect 35158 37816 35164 37828
rect 35216 37816 35222 37868
rect 37090 37816 37096 37868
rect 37148 37816 37154 37868
rect 37182 37816 37188 37868
rect 37240 37816 37246 37868
rect 37292 37856 37320 37896
rect 38930 37884 38936 37936
rect 38988 37884 38994 37936
rect 39942 37884 39948 37936
rect 40000 37924 40006 37936
rect 42153 37927 42211 37933
rect 40000 37896 40540 37924
rect 40000 37884 40006 37896
rect 37292 37828 40080 37856
rect 35342 37748 35348 37800
rect 35400 37748 35406 37800
rect 38746 37788 38752 37800
rect 38594 37760 38752 37788
rect 38746 37748 38752 37760
rect 38804 37748 38810 37800
rect 32784 37692 35572 37720
rect 31904 37680 31910 37692
rect 32125 37655 32183 37661
rect 32125 37652 32137 37655
rect 30484 37624 32137 37652
rect 30285 37615 30343 37621
rect 32125 37621 32137 37624
rect 32171 37621 32183 37655
rect 32125 37615 32183 37621
rect 33778 37612 33784 37664
rect 33836 37652 33842 37664
rect 34330 37652 34336 37664
rect 33836 37624 34336 37652
rect 33836 37612 33842 37624
rect 34330 37612 34336 37624
rect 34388 37612 34394 37664
rect 34514 37612 34520 37664
rect 34572 37652 34578 37664
rect 34609 37655 34667 37661
rect 34609 37652 34621 37655
rect 34572 37624 34621 37652
rect 34572 37612 34578 37624
rect 34609 37621 34621 37624
rect 34655 37621 34667 37655
rect 34609 37615 34667 37621
rect 34701 37655 34759 37661
rect 34701 37621 34713 37655
rect 34747 37652 34759 37655
rect 35434 37652 35440 37664
rect 34747 37624 35440 37652
rect 34747 37621 34759 37624
rect 34701 37615 34759 37621
rect 35434 37612 35440 37624
rect 35492 37612 35498 37664
rect 35544 37652 35572 37692
rect 37458 37680 37464 37732
rect 37516 37680 37522 37732
rect 39942 37652 39948 37664
rect 35544 37624 39948 37652
rect 39942 37612 39948 37624
rect 40000 37612 40006 37664
rect 40052 37652 40080 37828
rect 40402 37816 40408 37868
rect 40460 37816 40466 37868
rect 40512 37856 40540 37896
rect 42153 37893 42165 37927
rect 42199 37924 42211 37927
rect 42702 37924 42708 37936
rect 42199 37896 42708 37924
rect 42199 37893 42211 37896
rect 42153 37887 42211 37893
rect 41046 37856 41052 37868
rect 40512 37828 41052 37856
rect 41046 37816 41052 37828
rect 41104 37816 41110 37868
rect 41138 37816 41144 37868
rect 41196 37856 41202 37868
rect 41322 37856 41328 37868
rect 41196 37828 41328 37856
rect 41196 37816 41202 37828
rect 41322 37816 41328 37828
rect 41380 37856 41386 37868
rect 42168 37856 42196 37887
rect 42702 37884 42708 37896
rect 42760 37884 42766 37936
rect 44100 37924 44128 37964
rect 44174 37952 44180 38004
rect 44232 37952 44238 38004
rect 44450 37952 44456 38004
rect 44508 37952 44514 38004
rect 46385 37995 46443 38001
rect 46385 37961 46397 37995
rect 46431 37992 46443 37995
rect 46750 37992 46756 38004
rect 46431 37964 46756 37992
rect 46431 37961 46443 37964
rect 46385 37955 46443 37961
rect 46750 37952 46756 37964
rect 46808 37952 46814 38004
rect 49970 37992 49976 38004
rect 46860 37964 49976 37992
rect 46860 37924 46888 37964
rect 49970 37952 49976 37964
rect 50028 37952 50034 38004
rect 50144 37995 50202 38001
rect 50144 37961 50156 37995
rect 50190 37992 50202 37995
rect 50614 37992 50620 38004
rect 50190 37964 50620 37992
rect 50190 37961 50202 37964
rect 50144 37955 50202 37961
rect 50614 37952 50620 37964
rect 50672 37952 50678 38004
rect 50706 37952 50712 38004
rect 50764 37992 50770 38004
rect 51718 37992 51724 38004
rect 50764 37964 51724 37992
rect 50764 37952 50770 37964
rect 51718 37952 51724 37964
rect 51776 37952 51782 38004
rect 54386 37952 54392 38004
rect 54444 37952 54450 38004
rect 55769 37995 55827 38001
rect 55769 37961 55781 37995
rect 55815 37992 55827 37995
rect 56226 37992 56232 38004
rect 55815 37964 56232 37992
rect 55815 37961 55827 37964
rect 55769 37955 55827 37961
rect 56226 37952 56232 37964
rect 56284 37952 56290 38004
rect 57882 37952 57888 38004
rect 57940 37992 57946 38004
rect 63862 37992 63868 38004
rect 57940 37964 63868 37992
rect 57940 37952 57946 37964
rect 63862 37952 63868 37964
rect 63920 37952 63926 38004
rect 53834 37924 53840 37936
rect 44100 37896 46888 37924
rect 53668 37896 53840 37924
rect 41380 37828 42196 37856
rect 43625 37859 43683 37865
rect 41380 37816 41386 37828
rect 43625 37825 43637 37859
rect 43671 37856 43683 37859
rect 44082 37856 44088 37868
rect 43671 37828 44088 37856
rect 43671 37825 43683 37828
rect 43625 37819 43683 37825
rect 44082 37816 44088 37828
rect 44140 37816 44146 37868
rect 45002 37816 45008 37868
rect 45060 37816 45066 37868
rect 47118 37816 47124 37868
rect 47176 37856 47182 37868
rect 47854 37856 47860 37868
rect 47176 37828 47860 37856
rect 47176 37816 47182 37828
rect 47854 37816 47860 37828
rect 47912 37856 47918 37868
rect 48869 37859 48927 37865
rect 48869 37856 48881 37859
rect 47912 37828 48881 37856
rect 47912 37816 47918 37828
rect 48869 37825 48881 37828
rect 48915 37856 48927 37859
rect 49694 37856 49700 37868
rect 48915 37828 49700 37856
rect 48915 37825 48927 37828
rect 48869 37819 48927 37825
rect 49694 37816 49700 37828
rect 49752 37816 49758 37868
rect 50154 37856 50160 37868
rect 49804 37828 50160 37856
rect 42242 37748 42248 37800
rect 42300 37788 42306 37800
rect 43717 37791 43775 37797
rect 43717 37788 43729 37791
rect 42300 37760 43729 37788
rect 42300 37748 42306 37760
rect 43717 37757 43729 37760
rect 43763 37757 43775 37791
rect 43717 37751 43775 37757
rect 44818 37748 44824 37800
rect 44876 37748 44882 37800
rect 48133 37791 48191 37797
rect 48133 37757 48145 37791
rect 48179 37788 48191 37791
rect 49804 37788 49832 37828
rect 50154 37816 50160 37828
rect 50212 37816 50218 37868
rect 53668 37856 53696 37896
rect 53834 37884 53840 37896
rect 53892 37884 53898 37936
rect 56594 37924 56600 37936
rect 55140 37896 56600 37924
rect 52012 37828 53696 37856
rect 53745 37859 53803 37865
rect 48179 37760 49832 37788
rect 49881 37791 49939 37797
rect 48179 37757 48191 37760
rect 48133 37751 48191 37757
rect 49881 37757 49893 37791
rect 49927 37757 49939 37791
rect 49881 37751 49939 37757
rect 40681 37723 40739 37729
rect 40681 37689 40693 37723
rect 40727 37720 40739 37723
rect 40954 37720 40960 37732
rect 40727 37692 40960 37720
rect 40727 37689 40739 37692
rect 40681 37683 40739 37689
rect 40954 37680 40960 37692
rect 41012 37680 41018 37732
rect 41138 37680 41144 37732
rect 41196 37680 41202 37732
rect 44542 37680 44548 37732
rect 44600 37720 44606 37732
rect 44600 37692 46690 37720
rect 44600 37680 44606 37692
rect 47854 37680 47860 37732
rect 47912 37680 47918 37732
rect 48314 37680 48320 37732
rect 48372 37720 48378 37732
rect 49896 37720 49924 37751
rect 52012 37720 52040 37828
rect 53745 37825 53757 37859
rect 53791 37856 53803 37859
rect 54846 37856 54852 37868
rect 53791 37828 54852 37856
rect 53791 37825 53803 37828
rect 53745 37819 53803 37825
rect 54846 37816 54852 37828
rect 54904 37816 54910 37868
rect 55140 37865 55168 37896
rect 56594 37884 56600 37896
rect 56652 37884 56658 37936
rect 58434 37924 58440 37936
rect 57808 37896 58440 37924
rect 55125 37859 55183 37865
rect 55125 37825 55137 37859
rect 55171 37825 55183 37859
rect 57808 37856 57836 37896
rect 58434 37884 58440 37896
rect 58492 37884 58498 37936
rect 55125 37819 55183 37825
rect 55784 37828 57836 37856
rect 53466 37748 53472 37800
rect 53524 37788 53530 37800
rect 55214 37788 55220 37800
rect 53524 37760 55220 37788
rect 53524 37748 53530 37760
rect 55214 37748 55220 37760
rect 55272 37748 55278 37800
rect 48372 37692 49924 37720
rect 51382 37706 52040 37720
rect 51382 37692 52026 37706
rect 48372 37680 48378 37692
rect 53190 37680 53196 37732
rect 53248 37680 53254 37732
rect 53926 37680 53932 37732
rect 53984 37680 53990 37732
rect 54021 37723 54079 37729
rect 54021 37689 54033 37723
rect 54067 37720 54079 37723
rect 54202 37720 54208 37732
rect 54067 37692 54208 37720
rect 54067 37689 54079 37692
rect 54021 37683 54079 37689
rect 54202 37680 54208 37692
rect 54260 37680 54266 37732
rect 55122 37680 55128 37732
rect 55180 37720 55186 37732
rect 55309 37723 55367 37729
rect 55309 37720 55321 37723
rect 55180 37692 55321 37720
rect 55180 37680 55186 37692
rect 55309 37689 55321 37692
rect 55355 37689 55367 37723
rect 55309 37683 55367 37689
rect 55398 37680 55404 37732
rect 55456 37680 55462 37732
rect 42058 37652 42064 37664
rect 40052 37624 42064 37652
rect 42058 37612 42064 37624
rect 42116 37612 42122 37664
rect 43806 37612 43812 37664
rect 43864 37652 43870 37664
rect 44913 37655 44971 37661
rect 44913 37652 44925 37655
rect 43864 37624 44925 37652
rect 43864 37612 43870 37624
rect 44913 37621 44925 37624
rect 44959 37652 44971 37655
rect 45370 37652 45376 37664
rect 44959 37624 45376 37652
rect 44959 37621 44971 37624
rect 44913 37615 44971 37621
rect 45370 37612 45376 37624
rect 45428 37612 45434 37664
rect 47578 37612 47584 37664
rect 47636 37652 47642 37664
rect 48225 37655 48283 37661
rect 48225 37652 48237 37655
rect 47636 37624 48237 37652
rect 47636 37612 47642 37624
rect 48225 37621 48237 37624
rect 48271 37621 48283 37655
rect 48225 37615 48283 37621
rect 48406 37612 48412 37664
rect 48464 37652 48470 37664
rect 48593 37655 48651 37661
rect 48593 37652 48605 37655
rect 48464 37624 48605 37652
rect 48464 37612 48470 37624
rect 48593 37621 48605 37624
rect 48639 37621 48651 37655
rect 48593 37615 48651 37621
rect 48685 37655 48743 37661
rect 48685 37621 48697 37655
rect 48731 37652 48743 37655
rect 51629 37655 51687 37661
rect 51629 37652 51641 37655
rect 48731 37624 51641 37652
rect 48731 37621 48743 37624
rect 48685 37615 48743 37621
rect 51629 37621 51641 37624
rect 51675 37652 51687 37655
rect 51718 37652 51724 37664
rect 51675 37624 51724 37652
rect 51675 37621 51687 37624
rect 51629 37615 51687 37621
rect 51718 37612 51724 37624
rect 51776 37612 51782 37664
rect 51810 37612 51816 37664
rect 51868 37652 51874 37664
rect 55784 37652 55812 37828
rect 57882 37816 57888 37868
rect 57940 37816 57946 37868
rect 57974 37816 57980 37868
rect 58032 37856 58038 37868
rect 59725 37859 59783 37865
rect 59725 37856 59737 37859
rect 58032 37828 59737 37856
rect 58032 37816 58038 37828
rect 59725 37825 59737 37828
rect 59771 37856 59783 37859
rect 63126 37856 63132 37868
rect 59771 37828 63132 37856
rect 59771 37825 59783 37828
rect 59725 37819 59783 37825
rect 63126 37816 63132 37828
rect 63184 37816 63190 37868
rect 63678 37816 63684 37868
rect 63736 37816 63742 37868
rect 63770 37816 63776 37868
rect 63828 37816 63834 37868
rect 58342 37748 58348 37800
rect 58400 37748 58406 37800
rect 59909 37791 59967 37797
rect 59909 37757 59921 37791
rect 59955 37757 59967 37791
rect 59909 37751 59967 37757
rect 55858 37680 55864 37732
rect 55916 37680 55922 37732
rect 55950 37680 55956 37732
rect 56008 37720 56014 37732
rect 56008 37692 56442 37720
rect 56008 37680 56014 37692
rect 57330 37680 57336 37732
rect 57388 37720 57394 37732
rect 57609 37723 57667 37729
rect 57609 37720 57621 37723
rect 57388 37692 57621 37720
rect 57388 37680 57394 37692
rect 57609 37689 57621 37692
rect 57655 37689 57667 37723
rect 57609 37683 57667 37689
rect 59449 37723 59507 37729
rect 59449 37689 59461 37723
rect 59495 37720 59507 37723
rect 59814 37720 59820 37732
rect 59495 37692 59820 37720
rect 59495 37689 59507 37692
rect 59449 37683 59507 37689
rect 59814 37680 59820 37692
rect 59872 37680 59878 37732
rect 51868 37624 55812 37652
rect 55876 37652 55904 37680
rect 57790 37652 57796 37664
rect 55876 37624 57796 37652
rect 51868 37612 51874 37624
rect 57790 37612 57796 37624
rect 57848 37612 57854 37664
rect 57977 37655 58035 37661
rect 57977 37621 57989 37655
rect 58023 37652 58035 37655
rect 58526 37652 58532 37664
rect 58023 37624 58532 37652
rect 58023 37621 58035 37624
rect 57977 37615 58035 37621
rect 58526 37612 58532 37624
rect 58584 37652 58590 37664
rect 59924 37652 59952 37751
rect 59998 37748 60004 37800
rect 60056 37788 60062 37800
rect 66438 37788 66444 37800
rect 60056 37760 66444 37788
rect 60056 37748 60062 37760
rect 66438 37748 66444 37760
rect 66496 37748 66502 37800
rect 63865 37723 63923 37729
rect 63865 37689 63877 37723
rect 63911 37720 63923 37723
rect 65978 37720 65984 37732
rect 63911 37692 65984 37720
rect 63911 37689 63923 37692
rect 63865 37683 63923 37689
rect 65978 37680 65984 37692
rect 66036 37680 66042 37732
rect 58584 37624 59952 37652
rect 58584 37612 58590 37624
rect 60274 37612 60280 37664
rect 60332 37652 60338 37664
rect 60553 37655 60611 37661
rect 60553 37652 60565 37655
rect 60332 37624 60565 37652
rect 60332 37612 60338 37624
rect 60553 37621 60565 37624
rect 60599 37621 60611 37655
rect 60553 37615 60611 37621
rect 64230 37612 64236 37664
rect 64288 37612 64294 37664
rect 552 37562 66424 37584
rect 552 37510 2918 37562
rect 2970 37510 2982 37562
rect 3034 37510 3046 37562
rect 3098 37510 3110 37562
rect 3162 37510 3174 37562
rect 3226 37510 51918 37562
rect 51970 37510 51982 37562
rect 52034 37510 52046 37562
rect 52098 37510 52110 37562
rect 52162 37510 52174 37562
rect 52226 37510 65258 37562
rect 65310 37510 65322 37562
rect 65374 37510 65386 37562
rect 65438 37510 65450 37562
rect 65502 37510 65514 37562
rect 65566 37510 66424 37562
rect 552 37488 66424 37510
rect 9140 37420 12434 37448
rect 8754 37340 8760 37392
rect 8812 37340 8818 37392
rect 9030 37340 9036 37392
rect 9088 37380 9094 37392
rect 9140 37380 9168 37420
rect 12406 37380 12434 37420
rect 13538 37408 13544 37460
rect 13596 37448 13602 37460
rect 13596 37420 16620 37448
rect 13596 37408 13602 37420
rect 14274 37380 14280 37392
rect 9088 37352 9246 37380
rect 12406 37352 14280 37380
rect 9088 37340 9094 37352
rect 14274 37340 14280 37352
rect 14332 37340 14338 37392
rect 16592 37380 16620 37420
rect 17218 37408 17224 37460
rect 17276 37408 17282 37460
rect 17678 37408 17684 37460
rect 17736 37448 17742 37460
rect 18693 37451 18751 37457
rect 18693 37448 18705 37451
rect 17736 37420 18705 37448
rect 17736 37408 17742 37420
rect 18693 37417 18705 37420
rect 18739 37417 18751 37451
rect 18693 37411 18751 37417
rect 19061 37451 19119 37457
rect 19061 37417 19073 37451
rect 19107 37448 19119 37451
rect 19426 37448 19432 37460
rect 19107 37420 19432 37448
rect 19107 37417 19119 37420
rect 19061 37411 19119 37417
rect 17236 37380 17264 37408
rect 18138 37380 18144 37392
rect 16592 37352 17264 37380
rect 18078 37352 18144 37380
rect 8478 37272 8484 37324
rect 8536 37272 8542 37324
rect 10502 37272 10508 37324
rect 10560 37272 10566 37324
rect 13538 37272 13544 37324
rect 13596 37272 13602 37324
rect 16592 37321 16620 37352
rect 18138 37340 18144 37352
rect 18196 37340 18202 37392
rect 16577 37315 16635 37321
rect 16577 37281 16589 37315
rect 16623 37281 16635 37315
rect 19076 37312 19104 37411
rect 19426 37408 19432 37420
rect 19484 37408 19490 37460
rect 20622 37408 20628 37460
rect 20680 37448 20686 37460
rect 21453 37451 21511 37457
rect 21453 37448 21465 37451
rect 20680 37420 21465 37448
rect 20680 37408 20686 37420
rect 21453 37417 21465 37420
rect 21499 37417 21511 37451
rect 21453 37411 21511 37417
rect 21818 37408 21824 37460
rect 21876 37408 21882 37460
rect 23842 37408 23848 37460
rect 23900 37408 23906 37460
rect 24213 37451 24271 37457
rect 24213 37417 24225 37451
rect 24259 37448 24271 37451
rect 25130 37448 25136 37460
rect 24259 37420 25136 37448
rect 24259 37417 24271 37420
rect 24213 37411 24271 37417
rect 25130 37408 25136 37420
rect 25188 37408 25194 37460
rect 26510 37408 26516 37460
rect 26568 37448 26574 37460
rect 26881 37451 26939 37457
rect 26881 37448 26893 37451
rect 26568 37420 26893 37448
rect 26568 37408 26574 37420
rect 26881 37417 26893 37420
rect 26927 37417 26939 37451
rect 26881 37411 26939 37417
rect 27249 37451 27307 37457
rect 27249 37417 27261 37451
rect 27295 37448 27307 37451
rect 27798 37448 27804 37460
rect 27295 37420 27804 37448
rect 27295 37417 27307 37420
rect 27249 37411 27307 37417
rect 27798 37408 27804 37420
rect 27856 37408 27862 37460
rect 29178 37408 29184 37460
rect 29236 37448 29242 37460
rect 29914 37448 29920 37460
rect 29236 37420 29920 37448
rect 29236 37408 29242 37420
rect 29914 37408 29920 37420
rect 29972 37408 29978 37460
rect 31113 37451 31171 37457
rect 31113 37417 31125 37451
rect 31159 37417 31171 37451
rect 31113 37411 31171 37417
rect 31573 37451 31631 37457
rect 31573 37417 31585 37451
rect 31619 37448 31631 37451
rect 31662 37448 31668 37460
rect 31619 37420 31668 37448
rect 31619 37417 31631 37420
rect 31573 37411 31631 37417
rect 19153 37383 19211 37389
rect 19153 37349 19165 37383
rect 19199 37380 19211 37383
rect 19242 37380 19248 37392
rect 19199 37352 19248 37380
rect 19199 37349 19211 37352
rect 19153 37343 19211 37349
rect 19242 37340 19248 37352
rect 19300 37380 19306 37392
rect 21913 37383 21971 37389
rect 21913 37380 21925 37383
rect 19300 37352 21925 37380
rect 19300 37340 19306 37352
rect 21913 37349 21925 37352
rect 21959 37380 21971 37383
rect 28994 37380 29000 37392
rect 21959 37352 29000 37380
rect 21959 37349 21971 37352
rect 21913 37343 21971 37349
rect 28994 37340 29000 37352
rect 29052 37340 29058 37392
rect 16577 37275 16635 37281
rect 18340 37284 19104 37312
rect 13814 37204 13820 37256
rect 13872 37204 13878 37256
rect 15286 37204 15292 37256
rect 15344 37204 15350 37256
rect 16850 37204 16856 37256
rect 16908 37204 16914 37256
rect 18340 37253 18368 37284
rect 21818 37272 21824 37324
rect 21876 37312 21882 37324
rect 22278 37312 22284 37324
rect 21876 37284 22284 37312
rect 21876 37272 21882 37284
rect 22278 37272 22284 37284
rect 22336 37312 22342 37324
rect 24302 37312 24308 37324
rect 22336 37284 24308 37312
rect 22336 37272 22342 37284
rect 24302 37272 24308 37284
rect 24360 37272 24366 37324
rect 27341 37315 27399 37321
rect 27341 37281 27353 37315
rect 27387 37312 27399 37315
rect 27709 37315 27767 37321
rect 27709 37312 27721 37315
rect 27387 37284 27721 37312
rect 27387 37281 27399 37284
rect 27341 37275 27399 37281
rect 27709 37281 27721 37284
rect 27755 37281 27767 37315
rect 27709 37275 27767 37281
rect 28353 37315 28411 37321
rect 28353 37281 28365 37315
rect 28399 37312 28411 37315
rect 29196 37312 29224 37408
rect 29638 37340 29644 37392
rect 29696 37340 29702 37392
rect 30650 37340 30656 37392
rect 30708 37340 30714 37392
rect 28399 37284 29224 37312
rect 28399 37281 28411 37284
rect 28353 37275 28411 37281
rect 29362 37272 29368 37324
rect 29420 37272 29426 37324
rect 31128 37312 31156 37411
rect 31662 37408 31668 37420
rect 31720 37408 31726 37460
rect 31846 37408 31852 37460
rect 31904 37448 31910 37460
rect 31941 37451 31999 37457
rect 31941 37448 31953 37451
rect 31904 37420 31953 37448
rect 31904 37408 31910 37420
rect 31941 37417 31953 37420
rect 31987 37417 31999 37451
rect 31941 37411 31999 37417
rect 32033 37451 32091 37457
rect 32033 37417 32045 37451
rect 32079 37448 32091 37451
rect 32214 37448 32220 37460
rect 32079 37420 32220 37448
rect 32079 37417 32091 37420
rect 32033 37411 32091 37417
rect 32214 37408 32220 37420
rect 32272 37408 32278 37460
rect 32582 37408 32588 37460
rect 32640 37448 32646 37460
rect 34422 37448 34428 37460
rect 32640 37420 34428 37448
rect 32640 37408 32646 37420
rect 34422 37408 34428 37420
rect 34480 37408 34486 37460
rect 34514 37408 34520 37460
rect 34572 37408 34578 37460
rect 34885 37451 34943 37457
rect 34885 37417 34897 37451
rect 34931 37448 34943 37451
rect 35250 37448 35256 37460
rect 34931 37420 35256 37448
rect 34931 37417 34943 37420
rect 34885 37411 34943 37417
rect 35250 37408 35256 37420
rect 35308 37408 35314 37460
rect 35434 37408 35440 37460
rect 35492 37408 35498 37460
rect 35802 37408 35808 37460
rect 35860 37408 35866 37460
rect 36630 37408 36636 37460
rect 36688 37448 36694 37460
rect 38746 37448 38752 37460
rect 36688 37420 38752 37448
rect 36688 37408 36694 37420
rect 38746 37408 38752 37420
rect 38804 37408 38810 37460
rect 39114 37408 39120 37460
rect 39172 37448 39178 37460
rect 39301 37451 39359 37457
rect 39301 37448 39313 37451
rect 39172 37420 39313 37448
rect 39172 37408 39178 37420
rect 39301 37417 39313 37420
rect 39347 37417 39359 37451
rect 39301 37411 39359 37417
rect 40405 37451 40463 37457
rect 40405 37417 40417 37451
rect 40451 37448 40463 37451
rect 40770 37448 40776 37460
rect 40451 37420 40776 37448
rect 40451 37417 40463 37420
rect 40405 37411 40463 37417
rect 40770 37408 40776 37420
rect 40828 37408 40834 37460
rect 40865 37451 40923 37457
rect 40865 37417 40877 37451
rect 40911 37417 40923 37451
rect 40865 37411 40923 37417
rect 31754 37340 31760 37392
rect 31812 37380 31818 37392
rect 36725 37383 36783 37389
rect 36725 37380 36737 37383
rect 31812 37352 36737 37380
rect 31812 37340 31818 37352
rect 36725 37349 36737 37352
rect 36771 37349 36783 37383
rect 40497 37383 40555 37389
rect 40497 37380 40509 37383
rect 36725 37343 36783 37349
rect 36832 37352 40509 37380
rect 31846 37312 31852 37324
rect 31128 37284 31852 37312
rect 31846 37272 31852 37284
rect 31904 37272 31910 37324
rect 31938 37272 31944 37324
rect 31996 37312 32002 37324
rect 31996 37284 34376 37312
rect 31996 37272 32002 37284
rect 18325 37247 18383 37253
rect 18325 37213 18337 37247
rect 18371 37213 18383 37247
rect 18325 37207 18383 37213
rect 18874 37204 18880 37256
rect 18932 37244 18938 37256
rect 19245 37247 19303 37253
rect 19245 37244 19257 37247
rect 18932 37216 19257 37244
rect 18932 37204 18938 37216
rect 19245 37213 19257 37216
rect 19291 37213 19303 37247
rect 19245 37207 19303 37213
rect 20714 37204 20720 37256
rect 20772 37244 20778 37256
rect 21910 37244 21916 37256
rect 20772 37216 21916 37244
rect 20772 37204 20778 37216
rect 21910 37204 21916 37216
rect 21968 37244 21974 37256
rect 22005 37247 22063 37253
rect 22005 37244 22017 37247
rect 21968 37216 22017 37244
rect 21968 37204 21974 37216
rect 22005 37213 22017 37216
rect 22051 37213 22063 37247
rect 22005 37207 22063 37213
rect 24489 37247 24547 37253
rect 24489 37213 24501 37247
rect 24535 37244 24547 37247
rect 26234 37244 26240 37256
rect 24535 37216 26240 37244
rect 24535 37213 24547 37216
rect 24489 37207 24547 37213
rect 26234 37204 26240 37216
rect 26292 37204 26298 37256
rect 27430 37204 27436 37256
rect 27488 37204 27494 37256
rect 32030 37204 32036 37256
rect 32088 37244 32094 37256
rect 32125 37247 32183 37253
rect 32125 37244 32137 37247
rect 32088 37216 32137 37244
rect 32088 37204 32094 37216
rect 32125 37213 32137 37216
rect 32171 37213 32183 37247
rect 32125 37207 32183 37213
rect 34241 37247 34299 37253
rect 34241 37213 34253 37247
rect 34287 37213 34299 37247
rect 34241 37207 34299 37213
rect 33778 37176 33784 37188
rect 31404 37148 33784 37176
rect 27614 37068 27620 37120
rect 27672 37108 27678 37120
rect 31404 37108 31432 37148
rect 33778 37136 33784 37148
rect 33836 37136 33842 37188
rect 27672 37080 31432 37108
rect 27672 37068 27678 37080
rect 31478 37068 31484 37120
rect 31536 37108 31542 37120
rect 34256 37108 34284 37207
rect 34348 37176 34376 37284
rect 34514 37272 34520 37324
rect 34572 37312 34578 37324
rect 34977 37315 35035 37321
rect 34977 37312 34989 37315
rect 34572 37284 34989 37312
rect 34572 37272 34578 37284
rect 34977 37281 34989 37284
rect 35023 37281 35035 37315
rect 36832 37312 36860 37352
rect 40497 37349 40509 37352
rect 40543 37349 40555 37383
rect 40880 37380 40908 37411
rect 40954 37408 40960 37460
rect 41012 37408 41018 37460
rect 41417 37451 41475 37457
rect 41417 37448 41429 37451
rect 41156 37420 41429 37448
rect 41156 37380 41184 37420
rect 41417 37417 41429 37420
rect 41463 37417 41475 37451
rect 41417 37411 41475 37417
rect 46201 37451 46259 37457
rect 46201 37417 46213 37451
rect 46247 37448 46259 37451
rect 46247 37420 46520 37448
rect 46247 37417 46259 37420
rect 46201 37411 46259 37417
rect 46492 37380 46520 37420
rect 46566 37408 46572 37460
rect 46624 37448 46630 37460
rect 46661 37451 46719 37457
rect 46661 37448 46673 37451
rect 46624 37420 46673 37448
rect 46624 37408 46630 37420
rect 46661 37417 46673 37420
rect 46707 37417 46719 37451
rect 46661 37411 46719 37417
rect 47486 37408 47492 37460
rect 47544 37408 47550 37460
rect 47854 37408 47860 37460
rect 47912 37408 47918 37460
rect 50062 37408 50068 37460
rect 50120 37448 50126 37460
rect 50157 37451 50215 37457
rect 50157 37448 50169 37451
rect 50120 37420 50169 37448
rect 50120 37408 50126 37420
rect 50157 37417 50169 37420
rect 50203 37417 50215 37451
rect 50157 37411 50215 37417
rect 50617 37451 50675 37457
rect 50617 37417 50629 37451
rect 50663 37448 50675 37451
rect 50706 37448 50712 37460
rect 50663 37420 50712 37448
rect 50663 37417 50675 37420
rect 50617 37411 50675 37417
rect 50706 37408 50712 37420
rect 50764 37408 50770 37460
rect 50890 37408 50896 37460
rect 50948 37448 50954 37460
rect 51077 37451 51135 37457
rect 51077 37448 51089 37451
rect 50948 37420 51089 37448
rect 50948 37408 50954 37420
rect 51077 37417 51089 37420
rect 51123 37417 51135 37451
rect 51077 37411 51135 37417
rect 51537 37451 51595 37457
rect 51537 37417 51549 37451
rect 51583 37448 51595 37451
rect 53009 37451 53067 37457
rect 53009 37448 53021 37451
rect 51583 37420 53021 37448
rect 51583 37417 51595 37420
rect 51537 37411 51595 37417
rect 53009 37417 53021 37420
rect 53055 37417 53067 37451
rect 53009 37411 53067 37417
rect 53469 37451 53527 37457
rect 53469 37417 53481 37451
rect 53515 37448 53527 37451
rect 56778 37448 56784 37460
rect 53515 37420 56784 37448
rect 53515 37417 53527 37420
rect 53469 37411 53527 37417
rect 46750 37380 46756 37392
rect 40880 37352 41184 37380
rect 41248 37352 46428 37380
rect 46492 37352 46756 37380
rect 40497 37343 40555 37349
rect 34977 37275 35035 37281
rect 35084 37284 36860 37312
rect 34425 37247 34483 37253
rect 34425 37213 34437 37247
rect 34471 37244 34483 37247
rect 34698 37244 34704 37256
rect 34471 37216 34704 37244
rect 34471 37213 34483 37216
rect 34425 37207 34483 37213
rect 34698 37204 34704 37216
rect 34756 37204 34762 37256
rect 35084 37176 35112 37284
rect 36906 37272 36912 37324
rect 36964 37312 36970 37324
rect 36964 37284 38884 37312
rect 36964 37272 36970 37284
rect 35897 37247 35955 37253
rect 35897 37213 35909 37247
rect 35943 37213 35955 37247
rect 35897 37207 35955 37213
rect 34348 37148 35112 37176
rect 35345 37179 35403 37185
rect 35345 37145 35357 37179
rect 35391 37176 35403 37179
rect 35912 37176 35940 37207
rect 36078 37204 36084 37256
rect 36136 37204 36142 37256
rect 38473 37247 38531 37253
rect 38473 37213 38485 37247
rect 38519 37244 38531 37247
rect 38562 37244 38568 37256
rect 38519 37216 38568 37244
rect 38519 37213 38531 37216
rect 38473 37207 38531 37213
rect 38562 37204 38568 37216
rect 38620 37204 38626 37256
rect 38856 37244 38884 37284
rect 38930 37272 38936 37324
rect 38988 37312 38994 37324
rect 39669 37315 39727 37321
rect 39669 37312 39681 37315
rect 38988 37284 39681 37312
rect 38988 37272 38994 37284
rect 39669 37281 39681 37284
rect 39715 37281 39727 37315
rect 39669 37275 39727 37281
rect 39942 37272 39948 37324
rect 40000 37312 40006 37324
rect 41248 37312 41276 37352
rect 40000 37284 41276 37312
rect 40000 37272 40006 37284
rect 41322 37272 41328 37324
rect 41380 37272 41386 37324
rect 42058 37272 42064 37324
rect 42116 37312 42122 37324
rect 46293 37315 46351 37321
rect 46293 37312 46305 37315
rect 42116 37284 46305 37312
rect 42116 37272 42122 37284
rect 46293 37281 46305 37284
rect 46339 37281 46351 37315
rect 46400 37312 46428 37352
rect 46750 37340 46756 37352
rect 46808 37340 46814 37392
rect 47397 37383 47455 37389
rect 47397 37349 47409 37383
rect 47443 37380 47455 37383
rect 47578 37380 47584 37392
rect 47443 37352 47584 37380
rect 47443 37349 47455 37352
rect 47397 37343 47455 37349
rect 47578 37340 47584 37352
rect 47636 37340 47642 37392
rect 47688 37352 51074 37380
rect 47688 37312 47716 37352
rect 46400 37284 47716 37312
rect 46293 37275 46351 37281
rect 50062 37272 50068 37324
rect 50120 37312 50126 37324
rect 50709 37315 50767 37321
rect 50709 37312 50721 37315
rect 50120 37284 50721 37312
rect 50120 37272 50126 37284
rect 50709 37281 50721 37284
rect 50755 37281 50767 37315
rect 51046 37312 51074 37352
rect 51626 37340 51632 37392
rect 51684 37340 51690 37392
rect 51718 37340 51724 37392
rect 51776 37380 51782 37392
rect 52270 37380 52276 37392
rect 51776 37352 52276 37380
rect 51776 37340 51782 37352
rect 52270 37340 52276 37352
rect 52328 37380 52334 37392
rect 53377 37383 53435 37389
rect 53377 37380 53389 37383
rect 52328 37352 53389 37380
rect 52328 37340 52334 37352
rect 53377 37349 53389 37352
rect 53423 37349 53435 37383
rect 53377 37343 53435 37349
rect 51810 37312 51816 37324
rect 51046 37284 51816 37312
rect 50709 37275 50767 37281
rect 51810 37272 51816 37284
rect 51868 37272 51874 37324
rect 53190 37312 53196 37324
rect 52012 37284 53196 37312
rect 39761 37247 39819 37253
rect 39761 37244 39773 37247
rect 38856 37216 39773 37244
rect 39761 37213 39773 37216
rect 39807 37213 39819 37247
rect 39761 37207 39819 37213
rect 39853 37247 39911 37253
rect 39853 37213 39865 37247
rect 39899 37213 39911 37247
rect 39853 37207 39911 37213
rect 40313 37247 40371 37253
rect 40313 37213 40325 37247
rect 40359 37244 40371 37247
rect 40862 37244 40868 37256
rect 40359 37216 40868 37244
rect 40359 37213 40371 37216
rect 40313 37207 40371 37213
rect 39666 37176 39672 37188
rect 35391 37148 39672 37176
rect 35391 37145 35403 37148
rect 35345 37139 35403 37145
rect 39666 37136 39672 37148
rect 39724 37136 39730 37188
rect 34974 37108 34980 37120
rect 31536 37080 34980 37108
rect 31536 37068 31542 37080
rect 34974 37068 34980 37080
rect 35032 37108 35038 37120
rect 36078 37108 36084 37120
rect 35032 37080 36084 37108
rect 35032 37068 35038 37080
rect 36078 37068 36084 37080
rect 36136 37068 36142 37120
rect 36170 37068 36176 37120
rect 36228 37108 36234 37120
rect 39868 37108 39896 37207
rect 40862 37204 40868 37216
rect 40920 37204 40926 37256
rect 41230 37204 41236 37256
rect 41288 37244 41294 37256
rect 41509 37247 41567 37253
rect 41509 37244 41521 37247
rect 41288 37216 41521 37244
rect 41288 37204 41294 37216
rect 41509 37213 41521 37216
rect 41555 37213 41567 37247
rect 41509 37207 41567 37213
rect 46109 37247 46167 37253
rect 46109 37213 46121 37247
rect 46155 37244 46167 37247
rect 47118 37244 47124 37256
rect 46155 37216 47124 37244
rect 46155 37213 46167 37216
rect 46109 37207 46167 37213
rect 47118 37204 47124 37216
rect 47176 37204 47182 37256
rect 47302 37204 47308 37256
rect 47360 37204 47366 37256
rect 49694 37204 49700 37256
rect 49752 37244 49758 37256
rect 50522 37244 50528 37256
rect 49752 37216 50528 37244
rect 49752 37204 49758 37216
rect 50522 37204 50528 37216
rect 50580 37204 50586 37256
rect 51442 37204 51448 37256
rect 51500 37204 51506 37256
rect 40034 37136 40040 37188
rect 40092 37176 40098 37188
rect 52012 37185 52040 37284
rect 53190 37272 53196 37284
rect 53248 37272 53254 37324
rect 53484 37312 53512 37411
rect 56778 37408 56784 37420
rect 56836 37408 56842 37460
rect 57330 37408 57336 37460
rect 57388 37408 57394 37460
rect 57698 37408 57704 37460
rect 57756 37408 57762 37460
rect 57790 37408 57796 37460
rect 57848 37408 57854 37460
rect 58158 37408 58164 37460
rect 58216 37408 58222 37460
rect 58526 37408 58532 37460
rect 58584 37408 58590 37460
rect 58618 37408 58624 37460
rect 58676 37448 58682 37460
rect 59262 37448 59268 37460
rect 58676 37420 59268 37448
rect 58676 37408 58682 37420
rect 59262 37408 59268 37420
rect 59320 37448 59326 37460
rect 59357 37451 59415 37457
rect 59357 37448 59369 37451
rect 59320 37420 59369 37448
rect 59320 37408 59326 37420
rect 59357 37417 59369 37420
rect 59403 37417 59415 37451
rect 59357 37411 59415 37417
rect 59722 37408 59728 37460
rect 59780 37408 59786 37460
rect 59814 37408 59820 37460
rect 59872 37448 59878 37460
rect 59909 37451 59967 37457
rect 59909 37448 59921 37451
rect 59872 37420 59921 37448
rect 59872 37408 59878 37420
rect 59909 37417 59921 37420
rect 59955 37417 59967 37451
rect 59909 37411 59967 37417
rect 60274 37408 60280 37460
rect 60332 37408 60338 37460
rect 64877 37451 64935 37457
rect 64877 37417 64889 37451
rect 64923 37448 64935 37451
rect 65150 37448 65156 37460
rect 64923 37420 65156 37448
rect 64923 37417 64935 37420
rect 64877 37411 64935 37417
rect 65150 37408 65156 37420
rect 65208 37408 65214 37460
rect 55214 37380 55220 37392
rect 54496 37352 55220 37380
rect 53300 37284 53512 37312
rect 52917 37247 52975 37253
rect 52917 37213 52929 37247
rect 52963 37244 52975 37247
rect 53300 37244 53328 37284
rect 53650 37272 53656 37324
rect 53708 37312 53714 37324
rect 54496 37321 54524 37352
rect 55214 37340 55220 37352
rect 55272 37380 55278 37392
rect 56410 37380 56416 37392
rect 55272 37352 56416 37380
rect 55272 37340 55278 37352
rect 56410 37340 56416 37352
rect 56468 37340 56474 37392
rect 62758 37380 62764 37392
rect 56520 37352 62764 37380
rect 54481 37315 54539 37321
rect 53708 37284 54432 37312
rect 53708 37272 53714 37284
rect 52963 37216 53328 37244
rect 52963 37213 52975 37216
rect 52917 37207 52975 37213
rect 53558 37204 53564 37256
rect 53616 37204 53622 37256
rect 54404 37244 54432 37284
rect 54481 37281 54493 37315
rect 54527 37281 54539 37315
rect 54941 37315 54999 37321
rect 54941 37312 54953 37315
rect 54481 37275 54539 37281
rect 54588 37284 54953 37312
rect 54588 37244 54616 37284
rect 54941 37281 54953 37284
rect 54987 37312 54999 37315
rect 56520 37312 56548 37352
rect 62758 37340 62764 37352
rect 62816 37340 62822 37392
rect 64966 37380 64972 37392
rect 64630 37352 64972 37380
rect 64966 37340 64972 37352
rect 65024 37380 65030 37392
rect 65702 37380 65708 37392
rect 65024 37352 65708 37380
rect 65024 37340 65030 37352
rect 65702 37340 65708 37352
rect 65760 37340 65766 37392
rect 54987 37284 56548 37312
rect 54987 37281 54999 37284
rect 54941 37275 54999 37281
rect 57790 37272 57796 37324
rect 57848 37312 57854 37324
rect 59265 37315 59323 37321
rect 59265 37312 59277 37315
rect 57848 37284 59277 37312
rect 57848 37272 57854 37284
rect 59265 37281 59277 37284
rect 59311 37281 59323 37315
rect 59265 37275 59323 37281
rect 59906 37272 59912 37324
rect 59964 37312 59970 37324
rect 60369 37315 60427 37321
rect 60369 37312 60381 37315
rect 59964 37284 60381 37312
rect 59964 37272 59970 37284
rect 60369 37281 60381 37284
rect 60415 37281 60427 37315
rect 60369 37275 60427 37281
rect 63126 37272 63132 37324
rect 63184 37272 63190 37324
rect 65150 37272 65156 37324
rect 65208 37312 65214 37324
rect 65613 37315 65671 37321
rect 65613 37312 65625 37315
rect 65208 37284 65625 37312
rect 65208 37272 65214 37284
rect 65613 37281 65625 37284
rect 65659 37281 65671 37315
rect 65613 37275 65671 37281
rect 54404 37216 54616 37244
rect 54846 37204 54852 37256
rect 54904 37244 54910 37256
rect 57885 37247 57943 37253
rect 57885 37244 57897 37247
rect 54904 37216 57897 37244
rect 54904 37204 54910 37216
rect 57885 37213 57897 37216
rect 57931 37213 57943 37247
rect 57885 37207 57943 37213
rect 58710 37204 58716 37256
rect 58768 37204 58774 37256
rect 59081 37247 59139 37253
rect 59081 37213 59093 37247
rect 59127 37213 59139 37247
rect 59081 37207 59139 37213
rect 51997 37179 52055 37185
rect 40092 37148 51074 37176
rect 40092 37136 40098 37148
rect 36228 37080 39896 37108
rect 51046 37108 51074 37148
rect 51997 37145 52009 37179
rect 52043 37145 52055 37179
rect 51997 37139 52055 37145
rect 55876 37148 56548 37176
rect 55876 37108 55904 37148
rect 51046 37080 55904 37108
rect 36228 37068 36234 37080
rect 56410 37068 56416 37120
rect 56468 37068 56474 37120
rect 56520 37108 56548 37148
rect 56594 37136 56600 37188
rect 56652 37176 56658 37188
rect 57606 37176 57612 37188
rect 56652 37148 57612 37176
rect 56652 37136 56658 37148
rect 57606 37136 57612 37148
rect 57664 37176 57670 37188
rect 59096 37176 59124 37207
rect 60458 37204 60464 37256
rect 60516 37204 60522 37256
rect 63402 37204 63408 37256
rect 63460 37204 63466 37256
rect 59446 37176 59452 37188
rect 57664 37148 59452 37176
rect 57664 37136 57670 37148
rect 59446 37136 59452 37148
rect 59504 37176 59510 37188
rect 59504 37148 63080 37176
rect 59504 37136 59510 37148
rect 62942 37108 62948 37120
rect 56520 37080 62948 37108
rect 62942 37068 62948 37080
rect 63000 37068 63006 37120
rect 63052 37108 63080 37148
rect 64782 37108 64788 37120
rect 63052 37080 64788 37108
rect 64782 37068 64788 37080
rect 64840 37068 64846 37120
rect 64966 37068 64972 37120
rect 65024 37108 65030 37120
rect 65061 37111 65119 37117
rect 65061 37108 65073 37111
rect 65024 37080 65073 37108
rect 65024 37068 65030 37080
rect 65061 37077 65073 37080
rect 65107 37077 65119 37111
rect 65061 37071 65119 37077
rect 552 37018 66424 37040
rect 552 36966 1998 37018
rect 2050 36966 2062 37018
rect 2114 36966 2126 37018
rect 2178 36966 2190 37018
rect 2242 36966 2254 37018
rect 2306 36966 50998 37018
rect 51050 36966 51062 37018
rect 51114 36966 51126 37018
rect 51178 36966 51190 37018
rect 51242 36966 51254 37018
rect 51306 36966 64338 37018
rect 64390 36966 64402 37018
rect 64454 36966 64466 37018
rect 64518 36966 64530 37018
rect 64582 36966 64594 37018
rect 64646 36966 66424 37018
rect 552 36944 66424 36966
rect 10502 36864 10508 36916
rect 10560 36904 10566 36916
rect 24762 36904 24768 36916
rect 10560 36876 24768 36904
rect 10560 36864 10566 36876
rect 24762 36864 24768 36876
rect 24820 36864 24826 36916
rect 31662 36864 31668 36916
rect 31720 36904 31726 36916
rect 31938 36904 31944 36916
rect 31720 36876 31944 36904
rect 31720 36864 31726 36876
rect 31938 36864 31944 36876
rect 31996 36864 32002 36916
rect 51442 36864 51448 36916
rect 51500 36904 51506 36916
rect 54570 36904 54576 36916
rect 51500 36876 54576 36904
rect 51500 36864 51506 36876
rect 54570 36864 54576 36876
rect 54628 36864 54634 36916
rect 63402 36864 63408 36916
rect 63460 36904 63466 36916
rect 63865 36907 63923 36913
rect 63865 36904 63877 36907
rect 63460 36876 63877 36904
rect 63460 36864 63466 36876
rect 63865 36873 63877 36876
rect 63911 36873 63923 36907
rect 63865 36867 63923 36873
rect 25866 36796 25872 36848
rect 25924 36836 25930 36848
rect 35802 36836 35808 36848
rect 25924 36808 35808 36836
rect 25924 36796 25930 36808
rect 35802 36796 35808 36808
rect 35860 36796 35866 36848
rect 38654 36796 38660 36848
rect 38712 36836 38718 36848
rect 54588 36836 54616 36864
rect 60458 36836 60464 36848
rect 38712 36808 51074 36836
rect 54588 36808 60464 36836
rect 38712 36796 38718 36808
rect 19150 36728 19156 36780
rect 19208 36768 19214 36780
rect 38562 36768 38568 36780
rect 19208 36740 38568 36768
rect 19208 36728 19214 36740
rect 38562 36728 38568 36740
rect 38620 36728 38626 36780
rect 38746 36728 38752 36780
rect 38804 36768 38810 36780
rect 51046 36768 51074 36808
rect 60458 36796 60464 36808
rect 60516 36836 60522 36848
rect 60516 36808 64460 36836
rect 60516 36796 60522 36808
rect 63770 36768 63776 36780
rect 38804 36740 41414 36768
rect 51046 36740 63776 36768
rect 38804 36728 38810 36740
rect 14550 36660 14556 36712
rect 14608 36700 14614 36712
rect 38654 36700 38660 36712
rect 14608 36672 38660 36700
rect 14608 36660 14614 36672
rect 38654 36660 38660 36672
rect 38712 36660 38718 36712
rect 41386 36700 41414 36740
rect 63770 36728 63776 36740
rect 63828 36728 63834 36780
rect 64230 36728 64236 36780
rect 64288 36768 64294 36780
rect 64432 36777 64460 36808
rect 64782 36796 64788 36848
rect 64840 36836 64846 36848
rect 65886 36836 65892 36848
rect 64840 36808 65892 36836
rect 64840 36796 64846 36808
rect 65886 36796 65892 36808
rect 65944 36796 65950 36848
rect 64325 36771 64383 36777
rect 64325 36768 64337 36771
rect 64288 36740 64337 36768
rect 64288 36728 64294 36740
rect 64325 36737 64337 36740
rect 64371 36737 64383 36771
rect 64325 36731 64383 36737
rect 64417 36771 64475 36777
rect 64417 36737 64429 36771
rect 64463 36768 64475 36771
rect 64690 36768 64696 36780
rect 64463 36740 64696 36768
rect 64463 36737 64475 36740
rect 64417 36731 64475 36737
rect 64690 36728 64696 36740
rect 64748 36728 64754 36780
rect 65978 36728 65984 36780
rect 66036 36728 66042 36780
rect 41386 36672 65564 36700
rect 22002 36592 22008 36644
rect 22060 36632 22066 36644
rect 22060 36592 22094 36632
rect 30466 36592 30472 36644
rect 30524 36632 30530 36644
rect 34422 36632 34428 36644
rect 30524 36604 34428 36632
rect 30524 36592 30530 36604
rect 34422 36592 34428 36604
rect 34480 36592 34486 36644
rect 37642 36592 37648 36644
rect 37700 36632 37706 36644
rect 63494 36632 63500 36644
rect 37700 36604 63500 36632
rect 37700 36592 37706 36604
rect 63494 36592 63500 36604
rect 63552 36592 63558 36644
rect 64233 36635 64291 36641
rect 64233 36601 64245 36635
rect 64279 36632 64291 36635
rect 64966 36632 64972 36644
rect 64279 36604 64972 36632
rect 64279 36601 64291 36604
rect 64233 36595 64291 36601
rect 64966 36592 64972 36604
rect 65024 36592 65030 36644
rect 65536 36632 65564 36672
rect 66254 36632 66260 36644
rect 65536 36604 66260 36632
rect 66254 36592 66260 36604
rect 66312 36592 66318 36644
rect 22066 36428 22094 36592
rect 30282 36524 30288 36576
rect 30340 36564 30346 36576
rect 60826 36564 60832 36576
rect 30340 36536 60832 36564
rect 30340 36524 30346 36536
rect 60826 36524 60832 36536
rect 60884 36524 60890 36576
rect 65058 36524 65064 36576
rect 65116 36564 65122 36576
rect 65429 36567 65487 36573
rect 65429 36564 65441 36567
rect 65116 36536 65441 36564
rect 65116 36524 65122 36536
rect 65429 36533 65441 36536
rect 65475 36533 65487 36567
rect 65429 36527 65487 36533
rect 26970 36456 26976 36508
rect 27028 36496 27034 36508
rect 28810 36496 28816 36508
rect 27028 36468 28816 36496
rect 27028 36456 27034 36468
rect 28810 36456 28816 36468
rect 28868 36456 28874 36508
rect 30374 36456 30380 36508
rect 30432 36496 30438 36508
rect 37274 36496 37280 36508
rect 30432 36468 37280 36496
rect 30432 36456 30438 36468
rect 37274 36456 37280 36468
rect 37332 36456 37338 36508
rect 63572 36474 66424 36496
rect 33042 36428 33048 36440
rect 22066 36400 33048 36428
rect 33042 36388 33048 36400
rect 33100 36388 33106 36440
rect 63572 36422 65258 36474
rect 65310 36422 65322 36474
rect 65374 36422 65386 36474
rect 65438 36422 65450 36474
rect 65502 36422 65514 36474
rect 65566 36422 66424 36474
rect 63572 36400 66424 36422
rect 21634 36320 21640 36372
rect 21692 36360 21698 36372
rect 42702 36360 42708 36372
rect 21692 36332 42708 36360
rect 21692 36320 21698 36332
rect 42702 36320 42708 36332
rect 42760 36320 42766 36372
rect 65610 36320 65616 36372
rect 65668 36360 65674 36372
rect 65978 36360 65984 36372
rect 65668 36332 65984 36360
rect 65668 36320 65674 36332
rect 65978 36320 65984 36332
rect 66036 36320 66042 36372
rect 23198 36252 23204 36304
rect 23256 36292 23262 36304
rect 63586 36292 63592 36304
rect 23256 36264 63592 36292
rect 23256 36252 23262 36264
rect 63586 36252 63592 36264
rect 63644 36252 63650 36304
rect 65426 36292 65432 36304
rect 65366 36264 65432 36292
rect 65426 36252 65432 36264
rect 65484 36292 65490 36304
rect 65702 36292 65708 36304
rect 65484 36264 65708 36292
rect 65484 36252 65490 36264
rect 65702 36252 65708 36264
rect 65760 36252 65766 36304
rect 28718 36224 28724 36236
rect 22066 36196 28724 36224
rect 20070 35912 20076 35964
rect 20128 35952 20134 35964
rect 22066 35952 22094 36196
rect 28718 36184 28724 36196
rect 28776 36184 28782 36236
rect 28810 36184 28816 36236
rect 28868 36224 28874 36236
rect 33042 36224 33048 36236
rect 28868 36196 33048 36224
rect 28868 36184 28874 36196
rect 33042 36184 33048 36196
rect 33100 36184 33106 36236
rect 42610 36184 42616 36236
rect 42668 36224 42674 36236
rect 59354 36224 59360 36236
rect 42668 36196 59360 36224
rect 42668 36184 42674 36196
rect 59354 36184 59360 36196
rect 59412 36184 59418 36236
rect 23566 36116 23572 36168
rect 23624 36156 23630 36168
rect 62114 36156 62120 36168
rect 23624 36128 62120 36156
rect 23624 36116 23630 36128
rect 62114 36116 62120 36128
rect 62172 36116 62178 36168
rect 63862 36116 63868 36168
rect 63920 36116 63926 36168
rect 64141 36159 64199 36165
rect 64141 36125 64153 36159
rect 64187 36156 64199 36159
rect 64230 36156 64236 36168
rect 64187 36128 64236 36156
rect 64187 36125 64199 36128
rect 64141 36119 64199 36125
rect 64230 36116 64236 36128
rect 64288 36116 64294 36168
rect 24486 36048 24492 36100
rect 24544 36088 24550 36100
rect 63126 36088 63132 36100
rect 24544 36060 63132 36088
rect 24544 36048 24550 36060
rect 63126 36048 63132 36060
rect 63184 36048 63190 36100
rect 25222 35980 25228 36032
rect 25280 36020 25286 36032
rect 64782 36020 64788 36032
rect 25280 35992 64788 36020
rect 25280 35980 25286 35992
rect 64782 35980 64788 35992
rect 64840 35980 64846 36032
rect 20128 35924 22094 35952
rect 20128 35912 20134 35924
rect 24302 35912 24308 35964
rect 24360 35952 24366 35964
rect 24360 35924 30236 35952
rect 24360 35912 24366 35924
rect 21358 35844 21364 35896
rect 21416 35884 21422 35896
rect 21416 35856 22094 35884
rect 21416 35844 21422 35856
rect 22066 35816 22094 35856
rect 24762 35844 24768 35896
rect 24820 35884 24826 35896
rect 30098 35884 30104 35896
rect 24820 35856 30104 35884
rect 24820 35844 24826 35856
rect 30098 35844 30104 35856
rect 30156 35844 30162 35896
rect 30208 35884 30236 35924
rect 63572 35930 66424 35952
rect 36538 35884 36544 35896
rect 30208 35856 36544 35884
rect 36538 35844 36544 35856
rect 36596 35844 36602 35896
rect 63572 35878 64338 35930
rect 64390 35878 64402 35930
rect 64454 35878 64466 35930
rect 64518 35878 64530 35930
rect 64582 35878 64594 35930
rect 64646 35878 66424 35930
rect 63572 35856 66424 35878
rect 27614 35816 27620 35828
rect 22066 35788 27620 35816
rect 27614 35776 27620 35788
rect 27672 35776 27678 35828
rect 64230 35776 64236 35828
rect 64288 35816 64294 35828
rect 64693 35819 64751 35825
rect 64693 35816 64705 35819
rect 64288 35788 64705 35816
rect 64288 35776 64294 35788
rect 64693 35785 64705 35788
rect 64739 35785 64751 35819
rect 64693 35779 64751 35785
rect 8202 35708 8208 35760
rect 8260 35748 8266 35760
rect 14826 35748 14832 35760
rect 8260 35720 14832 35748
rect 8260 35708 8266 35720
rect 14826 35708 14832 35720
rect 14884 35708 14890 35760
rect 59354 35708 59360 35760
rect 59412 35748 59418 35760
rect 65702 35748 65708 35760
rect 59412 35720 65708 35748
rect 59412 35708 59418 35720
rect 65702 35708 65708 35720
rect 65760 35708 65766 35760
rect 22186 35640 22192 35692
rect 22244 35680 22250 35692
rect 42610 35680 42616 35692
rect 22244 35652 42616 35680
rect 22244 35640 22250 35652
rect 42610 35640 42616 35652
rect 42668 35640 42674 35692
rect 63678 35640 63684 35692
rect 63736 35680 63742 35692
rect 63957 35683 64015 35689
rect 63957 35680 63969 35683
rect 63736 35652 63969 35680
rect 63736 35640 63742 35652
rect 63957 35649 63969 35652
rect 64003 35649 64015 35683
rect 63957 35643 64015 35649
rect 64141 35683 64199 35689
rect 64141 35649 64153 35683
rect 64187 35680 64199 35683
rect 65150 35680 65156 35692
rect 64187 35652 65156 35680
rect 64187 35649 64199 35652
rect 64141 35643 64199 35649
rect 65150 35640 65156 35652
rect 65208 35640 65214 35692
rect 65337 35683 65395 35689
rect 65337 35649 65349 35683
rect 65383 35680 65395 35683
rect 65886 35680 65892 35692
rect 65383 35652 65892 35680
rect 65383 35649 65395 35652
rect 65337 35643 65395 35649
rect 65886 35640 65892 35652
rect 65944 35680 65950 35692
rect 66070 35680 66076 35692
rect 65944 35652 66076 35680
rect 65944 35640 65950 35652
rect 66070 35640 66076 35652
rect 66128 35640 66134 35692
rect 23014 35572 23020 35624
rect 23072 35612 23078 35624
rect 23072 35584 41414 35612
rect 23072 35572 23078 35584
rect 41386 35476 41414 35584
rect 62022 35572 62028 35624
rect 62080 35612 62086 35624
rect 64233 35615 64291 35621
rect 64233 35612 64245 35615
rect 62080 35584 64245 35612
rect 62080 35572 62086 35584
rect 64233 35581 64245 35584
rect 64279 35581 64291 35615
rect 64233 35575 64291 35581
rect 65058 35572 65064 35624
rect 65116 35572 65122 35624
rect 60826 35504 60832 35556
rect 60884 35544 60890 35556
rect 63494 35544 63500 35556
rect 60884 35516 63500 35544
rect 60884 35504 60890 35516
rect 63494 35504 63500 35516
rect 63552 35504 63558 35556
rect 65153 35547 65211 35553
rect 65153 35544 65165 35547
rect 64616 35516 65165 35544
rect 64230 35476 64236 35488
rect 41386 35448 64236 35476
rect 64230 35436 64236 35448
rect 64288 35436 64294 35488
rect 64616 35485 64644 35516
rect 65153 35513 65165 35516
rect 65199 35513 65211 35547
rect 65153 35507 65211 35513
rect 64601 35479 64659 35485
rect 64601 35445 64613 35479
rect 64647 35445 64659 35479
rect 64601 35439 64659 35445
rect 63572 35386 66424 35408
rect 63572 35334 65258 35386
rect 65310 35334 65322 35386
rect 65374 35334 65386 35386
rect 65438 35334 65450 35386
rect 65502 35334 65514 35386
rect 65566 35334 66424 35386
rect 63572 35312 66424 35334
rect 65794 35028 65800 35080
rect 65852 35068 65858 35080
rect 66070 35068 66076 35080
rect 65852 35040 66076 35068
rect 65852 35028 65858 35040
rect 66070 35028 66076 35040
rect 66128 35028 66134 35080
rect 62482 34892 62488 34944
rect 62540 34932 62546 34944
rect 64046 34932 64052 34944
rect 62540 34904 64052 34932
rect 62540 34892 62546 34904
rect 64046 34892 64052 34904
rect 64104 34892 64110 34944
rect 65610 34892 65616 34944
rect 65668 34932 65674 34944
rect 65794 34932 65800 34944
rect 65668 34904 65800 34932
rect 65668 34892 65674 34904
rect 65794 34892 65800 34904
rect 65852 34892 65858 34944
rect 63572 34842 66424 34864
rect 63572 34790 64338 34842
rect 64390 34790 64402 34842
rect 64454 34790 64466 34842
rect 64518 34790 64530 34842
rect 64582 34790 64594 34842
rect 64646 34790 66424 34842
rect 63572 34768 66424 34790
rect 63310 34688 63316 34740
rect 63368 34728 63374 34740
rect 65610 34728 65616 34740
rect 63368 34700 65616 34728
rect 63368 34688 63374 34700
rect 65610 34688 65616 34700
rect 65668 34688 65674 34740
rect 63862 34484 63868 34536
rect 63920 34484 63926 34536
rect 64138 34416 64144 34468
rect 64196 34416 64202 34468
rect 65150 34416 65156 34468
rect 65208 34416 65214 34468
rect 63572 34298 66424 34320
rect 63572 34246 65258 34298
rect 65310 34246 65322 34298
rect 65374 34246 65386 34298
rect 65438 34246 65450 34298
rect 65502 34246 65514 34298
rect 65566 34246 66424 34298
rect 63572 34224 66424 34246
rect 63957 34187 64015 34193
rect 63957 34153 63969 34187
rect 64003 34184 64015 34187
rect 64138 34184 64144 34196
rect 64003 34156 64144 34184
rect 64003 34153 64015 34156
rect 63957 34147 64015 34153
rect 64138 34144 64144 34156
rect 64196 34144 64202 34196
rect 64325 34051 64383 34057
rect 64325 34017 64337 34051
rect 64371 34048 64383 34051
rect 65061 34051 65119 34057
rect 65061 34048 65073 34051
rect 64371 34020 65073 34048
rect 64371 34017 64383 34020
rect 64325 34011 64383 34017
rect 65061 34017 65073 34020
rect 65107 34017 65119 34051
rect 65061 34011 65119 34017
rect 65610 34008 65616 34060
rect 65668 34008 65674 34060
rect 64417 33983 64475 33989
rect 64417 33949 64429 33983
rect 64463 33949 64475 33983
rect 64417 33943 64475 33949
rect 64601 33983 64659 33989
rect 64601 33949 64613 33983
rect 64647 33980 64659 33983
rect 64690 33980 64696 33992
rect 64647 33952 64696 33980
rect 64647 33949 64659 33952
rect 64601 33943 64659 33949
rect 64432 33844 64460 33943
rect 64690 33940 64696 33952
rect 64748 33940 64754 33992
rect 64690 33844 64696 33856
rect 64432 33816 64696 33844
rect 64690 33804 64696 33816
rect 64748 33804 64754 33856
rect 63572 33754 66424 33776
rect 63572 33702 64338 33754
rect 64390 33702 64402 33754
rect 64454 33702 64466 33754
rect 64518 33702 64530 33754
rect 64582 33702 64594 33754
rect 64646 33702 66424 33754
rect 63572 33680 66424 33702
rect 65978 33572 65984 33584
rect 64708 33544 65984 33572
rect 64708 33513 64736 33544
rect 65978 33532 65984 33544
rect 66036 33572 66042 33584
rect 66254 33572 66260 33584
rect 66036 33544 66260 33572
rect 66036 33532 66042 33544
rect 66254 33532 66260 33544
rect 66312 33532 66318 33584
rect 64693 33507 64751 33513
rect 64693 33473 64705 33507
rect 64739 33473 64751 33507
rect 64693 33467 64751 33473
rect 64782 33464 64788 33516
rect 64840 33504 64846 33516
rect 65058 33504 65064 33516
rect 64840 33476 65064 33504
rect 64840 33464 64846 33476
rect 65058 33464 65064 33476
rect 65116 33464 65122 33516
rect 64969 33439 65027 33445
rect 64969 33405 64981 33439
rect 65015 33436 65027 33439
rect 65610 33436 65616 33448
rect 65015 33408 65616 33436
rect 65015 33405 65027 33408
rect 64969 33399 65027 33405
rect 65610 33396 65616 33408
rect 65668 33396 65674 33448
rect 65978 33396 65984 33448
rect 66036 33396 66042 33448
rect 64877 33371 64935 33377
rect 64877 33337 64889 33371
rect 64923 33368 64935 33371
rect 66438 33368 66444 33380
rect 64923 33340 66444 33368
rect 64923 33337 64935 33340
rect 64877 33331 64935 33337
rect 66438 33328 66444 33340
rect 66496 33328 66502 33380
rect 65150 33260 65156 33312
rect 65208 33300 65214 33312
rect 65337 33303 65395 33309
rect 65337 33300 65349 33303
rect 65208 33272 65349 33300
rect 65208 33260 65214 33272
rect 65337 33269 65349 33272
rect 65383 33269 65395 33303
rect 65337 33263 65395 33269
rect 65429 33303 65487 33309
rect 65429 33269 65441 33303
rect 65475 33300 65487 33303
rect 65610 33300 65616 33312
rect 65475 33272 65616 33300
rect 65475 33269 65487 33272
rect 65429 33263 65487 33269
rect 65610 33260 65616 33272
rect 65668 33260 65674 33312
rect 62850 33192 62856 33244
rect 62908 33232 62914 33244
rect 63402 33232 63408 33244
rect 62908 33204 63408 33232
rect 62908 33192 62914 33204
rect 63402 33192 63408 33204
rect 63460 33192 63466 33244
rect 63572 33210 66424 33232
rect 63572 33158 65258 33210
rect 65310 33158 65322 33210
rect 65374 33158 65386 33210
rect 65438 33158 65450 33210
rect 65502 33158 65514 33210
rect 65566 33158 66424 33210
rect 63572 33136 66424 33158
rect 66070 33028 66076 33040
rect 65458 33000 66076 33028
rect 66070 32988 66076 33000
rect 66128 32988 66134 33040
rect 63954 32852 63960 32904
rect 64012 32852 64018 32904
rect 64233 32895 64291 32901
rect 64233 32861 64245 32895
rect 64279 32892 64291 32895
rect 64874 32892 64880 32904
rect 64279 32864 64880 32892
rect 64279 32861 64291 32864
rect 64233 32855 64291 32861
rect 64874 32852 64880 32864
rect 64932 32852 64938 32904
rect 65242 32716 65248 32768
rect 65300 32756 65306 32768
rect 65705 32759 65763 32765
rect 65705 32756 65717 32759
rect 65300 32728 65717 32756
rect 65300 32716 65306 32728
rect 65705 32725 65717 32728
rect 65751 32756 65763 32759
rect 65978 32756 65984 32768
rect 65751 32728 65984 32756
rect 65751 32725 65763 32728
rect 65705 32719 65763 32725
rect 65978 32716 65984 32728
rect 66036 32716 66042 32768
rect 63572 32666 66424 32688
rect 63572 32614 64338 32666
rect 64390 32614 64402 32666
rect 64454 32614 64466 32666
rect 64518 32614 64530 32666
rect 64582 32614 64594 32666
rect 64646 32614 66424 32666
rect 63572 32592 66424 32614
rect 64690 32512 64696 32564
rect 64748 32512 64754 32564
rect 64874 32512 64880 32564
rect 64932 32552 64938 32564
rect 64969 32555 65027 32561
rect 64969 32552 64981 32555
rect 64932 32524 64981 32552
rect 64932 32512 64938 32524
rect 64969 32521 64981 32524
rect 65015 32521 65027 32555
rect 64969 32515 65027 32521
rect 65978 32484 65984 32496
rect 64156 32456 65984 32484
rect 64156 32425 64184 32456
rect 65978 32444 65984 32456
rect 66036 32484 66042 32496
rect 66254 32484 66260 32496
rect 66036 32456 66260 32484
rect 66036 32444 66042 32456
rect 66254 32444 66260 32456
rect 66312 32444 66318 32496
rect 64141 32419 64199 32425
rect 64141 32385 64153 32419
rect 64187 32385 64199 32419
rect 64141 32379 64199 32385
rect 65150 32376 65156 32428
rect 65208 32416 65214 32428
rect 65429 32419 65487 32425
rect 65429 32416 65441 32419
rect 65208 32388 65441 32416
rect 65208 32376 65214 32388
rect 65429 32385 65441 32388
rect 65475 32385 65487 32419
rect 65429 32379 65487 32385
rect 65521 32419 65579 32425
rect 65521 32385 65533 32419
rect 65567 32416 65579 32419
rect 65886 32416 65892 32428
rect 65567 32388 65892 32416
rect 65567 32385 65579 32388
rect 65521 32379 65579 32385
rect 64233 32351 64291 32357
rect 64233 32317 64245 32351
rect 64279 32348 64291 32351
rect 65242 32348 65248 32360
rect 64279 32320 65248 32348
rect 64279 32317 64291 32320
rect 64233 32311 64291 32317
rect 65242 32308 65248 32320
rect 65300 32308 65306 32360
rect 65337 32351 65395 32357
rect 65337 32317 65349 32351
rect 65383 32348 65395 32351
rect 65610 32348 65616 32360
rect 65383 32320 65616 32348
rect 65383 32317 65395 32320
rect 65337 32311 65395 32317
rect 65610 32308 65616 32320
rect 65668 32308 65674 32360
rect 64325 32283 64383 32289
rect 64325 32249 64337 32283
rect 64371 32280 64383 32283
rect 64785 32283 64843 32289
rect 64785 32280 64797 32283
rect 64371 32252 64797 32280
rect 64371 32249 64383 32252
rect 64325 32243 64383 32249
rect 64785 32249 64797 32252
rect 64831 32280 64843 32283
rect 64874 32280 64880 32292
rect 64831 32252 64880 32280
rect 64831 32249 64843 32252
rect 64785 32243 64843 32249
rect 64874 32240 64880 32252
rect 64932 32280 64938 32292
rect 65702 32280 65708 32292
rect 64932 32252 65708 32280
rect 64932 32240 64938 32252
rect 65702 32240 65708 32252
rect 65760 32240 65766 32292
rect 65610 32172 65616 32224
rect 65668 32212 65674 32224
rect 65812 32212 65840 32388
rect 65886 32376 65892 32388
rect 65944 32376 65950 32428
rect 65668 32184 65840 32212
rect 65668 32172 65674 32184
rect 63572 32122 66424 32144
rect 63572 32070 65258 32122
rect 65310 32070 65322 32122
rect 65374 32070 65386 32122
rect 65438 32070 65450 32122
rect 65502 32070 65514 32122
rect 65566 32070 66424 32122
rect 63572 32048 66424 32070
rect 63862 31968 63868 32020
rect 63920 32008 63926 32020
rect 64046 32008 64052 32020
rect 63920 31980 64052 32008
rect 63920 31968 63926 31980
rect 64046 31968 64052 31980
rect 64104 32008 64110 32020
rect 65429 32011 65487 32017
rect 65429 32008 65441 32011
rect 64104 31980 65441 32008
rect 64104 31968 64110 31980
rect 65429 31977 65441 31980
rect 65475 31977 65487 32011
rect 65429 31971 65487 31977
rect 64141 31943 64199 31949
rect 64141 31909 64153 31943
rect 64187 31940 64199 31943
rect 64966 31940 64972 31952
rect 64187 31912 64972 31940
rect 64187 31909 64199 31912
rect 64141 31903 64199 31909
rect 64966 31900 64972 31912
rect 65024 31900 65030 31952
rect 63678 31832 63684 31884
rect 63736 31872 63742 31884
rect 63862 31872 63868 31884
rect 63736 31844 63868 31872
rect 63736 31832 63742 31844
rect 63862 31832 63868 31844
rect 63920 31832 63926 31884
rect 64049 31875 64107 31881
rect 64049 31841 64061 31875
rect 64095 31872 64107 31875
rect 64874 31872 64880 31884
rect 64095 31844 64880 31872
rect 64095 31841 64107 31844
rect 64049 31835 64107 31841
rect 64874 31832 64880 31844
rect 64932 31832 64938 31884
rect 63572 31578 66424 31600
rect 63572 31526 64338 31578
rect 64390 31526 64402 31578
rect 64454 31526 64466 31578
rect 64518 31526 64530 31578
rect 64582 31526 64594 31578
rect 64646 31526 66424 31578
rect 63572 31504 66424 31526
rect 64601 31399 64659 31405
rect 64601 31365 64613 31399
rect 64647 31396 64659 31399
rect 65058 31396 65064 31408
rect 64647 31368 65064 31396
rect 64647 31365 64659 31368
rect 64601 31359 64659 31365
rect 65058 31356 65064 31368
rect 65116 31356 65122 31408
rect 64874 31288 64880 31340
rect 64932 31328 64938 31340
rect 65245 31331 65303 31337
rect 65245 31328 65257 31331
rect 64932 31300 65257 31328
rect 64932 31288 64938 31300
rect 65245 31297 65257 31300
rect 65291 31328 65303 31331
rect 65978 31328 65984 31340
rect 65291 31300 65984 31328
rect 65291 31297 65303 31300
rect 65245 31291 65303 31297
rect 65978 31288 65984 31300
rect 66036 31288 66042 31340
rect 66070 31288 66076 31340
rect 66128 31288 66134 31340
rect 65061 31263 65119 31269
rect 65061 31229 65073 31263
rect 65107 31260 65119 31263
rect 65794 31260 65800 31272
rect 65107 31232 65800 31260
rect 65107 31229 65119 31232
rect 65061 31223 65119 31229
rect 65794 31220 65800 31232
rect 65852 31220 65858 31272
rect 64969 31195 65027 31201
rect 64969 31161 64981 31195
rect 65015 31192 65027 31195
rect 65702 31192 65708 31204
rect 65015 31164 65708 31192
rect 65015 31161 65027 31164
rect 64969 31155 65027 31161
rect 65702 31152 65708 31164
rect 65760 31152 65766 31204
rect 65794 31084 65800 31136
rect 65852 31124 65858 31136
rect 66088 31124 66116 31288
rect 65852 31096 66116 31124
rect 65852 31084 65858 31096
rect 63572 31034 66424 31056
rect 62574 30948 62580 31000
rect 62632 30988 62638 31000
rect 63218 30988 63224 31000
rect 62632 30960 63224 30988
rect 62632 30948 62638 30960
rect 63218 30948 63224 30960
rect 63276 30948 63282 31000
rect 63572 30982 65258 31034
rect 65310 30982 65322 31034
rect 65374 30982 65386 31034
rect 65438 30982 65450 31034
rect 65502 30982 65514 31034
rect 65566 30982 66424 31034
rect 63572 30960 66424 30982
rect 65794 30852 65800 30864
rect 65550 30824 65800 30852
rect 65794 30812 65800 30824
rect 65852 30812 65858 30864
rect 63954 30744 63960 30796
rect 64012 30784 64018 30796
rect 64049 30787 64107 30793
rect 64049 30784 64061 30787
rect 64012 30756 64061 30784
rect 64012 30744 64018 30756
rect 64049 30753 64061 30756
rect 64095 30753 64107 30787
rect 64049 30747 64107 30753
rect 64325 30719 64383 30725
rect 64325 30685 64337 30719
rect 64371 30716 64383 30719
rect 64690 30716 64696 30728
rect 64371 30688 64696 30716
rect 64371 30685 64383 30688
rect 64325 30679 64383 30685
rect 64690 30676 64696 30688
rect 64748 30676 64754 30728
rect 65797 30583 65855 30589
rect 65797 30549 65809 30583
rect 65843 30580 65855 30583
rect 65978 30580 65984 30592
rect 65843 30552 65984 30580
rect 65843 30549 65855 30552
rect 65797 30543 65855 30549
rect 65978 30540 65984 30552
rect 66036 30540 66042 30592
rect 63572 30490 66424 30512
rect 63572 30438 64338 30490
rect 64390 30438 64402 30490
rect 64454 30438 64466 30490
rect 64518 30438 64530 30490
rect 64582 30438 64594 30490
rect 64646 30438 66424 30490
rect 63572 30416 66424 30438
rect 64601 30379 64659 30385
rect 64601 30345 64613 30379
rect 64647 30376 64659 30379
rect 64690 30376 64696 30388
rect 64647 30348 64696 30376
rect 64647 30345 64659 30348
rect 64601 30339 64659 30345
rect 64690 30336 64696 30348
rect 64748 30336 64754 30388
rect 65058 30200 65064 30252
rect 65116 30200 65122 30252
rect 65245 30243 65303 30249
rect 65245 30209 65257 30243
rect 65291 30240 65303 30243
rect 65610 30240 65616 30252
rect 65291 30212 65616 30240
rect 65291 30209 65303 30212
rect 65245 30203 65303 30209
rect 65610 30200 65616 30212
rect 65668 30200 65674 30252
rect 65978 30132 65984 30184
rect 66036 30132 66042 30184
rect 64969 30107 65027 30113
rect 64969 30073 64981 30107
rect 65015 30104 65027 30107
rect 65429 30107 65487 30113
rect 65429 30104 65441 30107
rect 65015 30076 65441 30104
rect 65015 30073 65027 30076
rect 64969 30067 65027 30073
rect 65429 30073 65441 30076
rect 65475 30073 65487 30107
rect 65429 30067 65487 30073
rect 63572 29946 66424 29968
rect 63572 29894 65258 29946
rect 65310 29894 65322 29946
rect 65374 29894 65386 29946
rect 65438 29894 65450 29946
rect 65502 29894 65514 29946
rect 65566 29894 66424 29946
rect 63572 29872 66424 29894
rect 64969 29767 65027 29773
rect 64969 29733 64981 29767
rect 65015 29764 65027 29767
rect 65058 29764 65064 29776
rect 65015 29736 65064 29764
rect 65015 29733 65027 29736
rect 64969 29727 65027 29733
rect 65058 29724 65064 29736
rect 65116 29724 65122 29776
rect 64877 29699 64935 29705
rect 64877 29665 64889 29699
rect 64923 29696 64935 29699
rect 65429 29699 65487 29705
rect 65429 29696 65441 29699
rect 64923 29668 65441 29696
rect 64923 29665 64935 29668
rect 64877 29659 64935 29665
rect 65429 29665 65441 29668
rect 65475 29665 65487 29699
rect 65429 29659 65487 29665
rect 65153 29631 65211 29637
rect 65153 29597 65165 29631
rect 65199 29628 65211 29631
rect 65610 29628 65616 29640
rect 65199 29600 65616 29628
rect 65199 29597 65211 29600
rect 65153 29591 65211 29597
rect 65610 29588 65616 29600
rect 65668 29588 65674 29640
rect 65702 29588 65708 29640
rect 65760 29628 65766 29640
rect 65981 29631 66039 29637
rect 65981 29628 65993 29631
rect 65760 29600 65993 29628
rect 65760 29588 65766 29600
rect 65981 29597 65993 29600
rect 66027 29597 66039 29631
rect 65981 29591 66039 29597
rect 64509 29495 64567 29501
rect 64509 29461 64521 29495
rect 64555 29492 64567 29495
rect 64690 29492 64696 29504
rect 64555 29464 64696 29492
rect 64555 29461 64567 29464
rect 64509 29455 64567 29461
rect 64690 29452 64696 29464
rect 64748 29452 64754 29504
rect 63572 29402 66424 29424
rect 63572 29350 64338 29402
rect 64390 29350 64402 29402
rect 64454 29350 64466 29402
rect 64518 29350 64530 29402
rect 64582 29350 64594 29402
rect 64646 29350 66424 29402
rect 63572 29328 66424 29350
rect 64046 29112 64052 29164
rect 64104 29112 64110 29164
rect 64325 29155 64383 29161
rect 64325 29121 64337 29155
rect 64371 29152 64383 29155
rect 64690 29152 64696 29164
rect 64371 29124 64696 29152
rect 64371 29121 64383 29124
rect 64325 29115 64383 29121
rect 64690 29112 64696 29124
rect 64748 29112 64754 29164
rect 65702 29112 65708 29164
rect 65760 29152 65766 29164
rect 65797 29155 65855 29161
rect 65797 29152 65809 29155
rect 65760 29124 65809 29152
rect 65760 29112 65766 29124
rect 65797 29121 65809 29124
rect 65843 29121 65855 29155
rect 65797 29115 65855 29121
rect 65794 29016 65800 29028
rect 65550 28988 65800 29016
rect 65794 28976 65800 28988
rect 65852 29016 65858 29028
rect 66162 29016 66168 29028
rect 65852 28988 66168 29016
rect 65852 28976 65858 28988
rect 66162 28976 66168 28988
rect 66220 28976 66226 29028
rect 63572 28858 66424 28880
rect 63572 28806 65258 28858
rect 65310 28806 65322 28858
rect 65374 28806 65386 28858
rect 65438 28806 65450 28858
rect 65502 28806 65514 28858
rect 65566 28806 66424 28858
rect 63572 28784 66424 28806
rect 65058 28704 65064 28756
rect 65116 28704 65122 28756
rect 64693 28679 64751 28685
rect 64693 28645 64705 28679
rect 64739 28676 64751 28679
rect 65150 28676 65156 28688
rect 64739 28648 65156 28676
rect 64739 28645 64751 28648
rect 64693 28639 64751 28645
rect 65150 28636 65156 28648
rect 65208 28636 65214 28688
rect 64601 28611 64659 28617
rect 64601 28577 64613 28611
rect 64647 28608 64659 28611
rect 65978 28608 65984 28620
rect 64647 28580 65984 28608
rect 64647 28577 64659 28580
rect 64601 28571 64659 28577
rect 65978 28568 65984 28580
rect 66036 28568 66042 28620
rect 64509 28543 64567 28549
rect 64509 28509 64521 28543
rect 64555 28509 64567 28543
rect 64509 28503 64567 28509
rect 64524 28472 64552 28503
rect 64966 28472 64972 28484
rect 64524 28444 64972 28472
rect 64966 28432 64972 28444
rect 65024 28432 65030 28484
rect 63572 28314 66424 28336
rect 63572 28262 64338 28314
rect 64390 28262 64402 28314
rect 64454 28262 64466 28314
rect 64518 28262 64530 28314
rect 64582 28262 64594 28314
rect 64646 28262 66424 28314
rect 63572 28240 66424 28262
rect 63572 27770 66424 27792
rect 63572 27718 65258 27770
rect 65310 27718 65322 27770
rect 65374 27718 65386 27770
rect 65438 27718 65450 27770
rect 65502 27718 65514 27770
rect 65566 27718 66424 27770
rect 63572 27696 66424 27718
rect 62850 27548 62856 27600
rect 62908 27588 62914 27600
rect 63494 27588 63500 27600
rect 62908 27560 63500 27588
rect 62908 27548 62914 27560
rect 63494 27548 63500 27560
rect 63552 27548 63558 27600
rect 63572 27226 66424 27248
rect 63572 27174 64338 27226
rect 64390 27174 64402 27226
rect 64454 27174 64466 27226
rect 64518 27174 64530 27226
rect 64582 27174 64594 27226
rect 64646 27174 66424 27226
rect 63572 27152 66424 27174
rect 64601 27047 64659 27053
rect 64601 27013 64613 27047
rect 64647 27044 64659 27047
rect 65058 27044 65064 27056
rect 64647 27016 65064 27044
rect 64647 27013 64659 27016
rect 64601 27007 64659 27013
rect 65058 27004 65064 27016
rect 65116 27004 65122 27056
rect 64966 26936 64972 26988
rect 65024 26976 65030 26988
rect 65153 26979 65211 26985
rect 65153 26976 65165 26979
rect 65024 26948 65165 26976
rect 65024 26936 65030 26948
rect 65153 26945 65165 26948
rect 65199 26945 65211 26979
rect 65153 26939 65211 26945
rect 65061 26911 65119 26917
rect 65061 26877 65073 26911
rect 65107 26908 65119 26911
rect 65702 26908 65708 26920
rect 65107 26880 65708 26908
rect 65107 26877 65119 26880
rect 65061 26871 65119 26877
rect 65702 26868 65708 26880
rect 65760 26868 65766 26920
rect 64969 26843 65027 26849
rect 64969 26809 64981 26843
rect 65015 26840 65027 26843
rect 65794 26840 65800 26852
rect 65015 26812 65800 26840
rect 65015 26809 65027 26812
rect 64969 26803 65027 26809
rect 65794 26800 65800 26812
rect 65852 26800 65858 26852
rect 63572 26682 66424 26704
rect 63572 26630 65258 26682
rect 65310 26630 65322 26682
rect 65374 26630 65386 26682
rect 65438 26630 65450 26682
rect 65502 26630 65514 26682
rect 65566 26630 66424 26682
rect 63572 26608 66424 26630
rect 64966 26528 64972 26580
rect 65024 26568 65030 26580
rect 65610 26568 65616 26580
rect 65024 26540 65616 26568
rect 65024 26528 65030 26540
rect 65610 26528 65616 26540
rect 65668 26528 65674 26580
rect 66162 26500 66168 26512
rect 65550 26486 66168 26500
rect 65536 26472 66168 26486
rect 64046 26324 64052 26376
rect 64104 26324 64110 26376
rect 64325 26367 64383 26373
rect 64325 26333 64337 26367
rect 64371 26364 64383 26367
rect 64690 26364 64696 26376
rect 64371 26336 64696 26364
rect 64371 26333 64383 26336
rect 64325 26327 64383 26333
rect 64690 26324 64696 26336
rect 64748 26324 64754 26376
rect 64966 26324 64972 26376
rect 65024 26364 65030 26376
rect 65536 26364 65564 26472
rect 66162 26460 66168 26472
rect 66220 26460 66226 26512
rect 65024 26336 65564 26364
rect 65024 26324 65030 26336
rect 65797 26231 65855 26237
rect 65797 26197 65809 26231
rect 65843 26228 65855 26231
rect 65978 26228 65984 26240
rect 65843 26200 65984 26228
rect 65843 26197 65855 26200
rect 65797 26191 65855 26197
rect 65978 26188 65984 26200
rect 66036 26188 66042 26240
rect 63572 26138 66424 26160
rect 63572 26086 64338 26138
rect 64390 26086 64402 26138
rect 64454 26086 64466 26138
rect 64518 26086 64530 26138
rect 64582 26086 64594 26138
rect 64646 26086 66424 26138
rect 63572 26064 66424 26086
rect 64601 26027 64659 26033
rect 64601 25993 64613 26027
rect 64647 26024 64659 26027
rect 64690 26024 64696 26036
rect 64647 25996 64696 26024
rect 64647 25993 64659 25996
rect 64601 25987 64659 25993
rect 64690 25984 64696 25996
rect 64748 25984 64754 26036
rect 65058 25848 65064 25900
rect 65116 25848 65122 25900
rect 65150 25848 65156 25900
rect 65208 25888 65214 25900
rect 65245 25891 65303 25897
rect 65245 25888 65257 25891
rect 65208 25860 65257 25888
rect 65208 25848 65214 25860
rect 65245 25857 65257 25860
rect 65291 25888 65303 25891
rect 65702 25888 65708 25900
rect 65291 25860 65708 25888
rect 65291 25857 65303 25860
rect 65245 25851 65303 25857
rect 65702 25848 65708 25860
rect 65760 25848 65766 25900
rect 65978 25780 65984 25832
rect 66036 25780 66042 25832
rect 64969 25687 65027 25693
rect 64969 25653 64981 25687
rect 65015 25684 65027 25687
rect 65429 25687 65487 25693
rect 65429 25684 65441 25687
rect 65015 25656 65441 25684
rect 65015 25653 65027 25656
rect 64969 25647 65027 25653
rect 65429 25653 65441 25656
rect 65475 25653 65487 25687
rect 65429 25647 65487 25653
rect 63572 25594 66424 25616
rect 63572 25542 65258 25594
rect 65310 25542 65322 25594
rect 65374 25542 65386 25594
rect 65438 25542 65450 25594
rect 65502 25542 65514 25594
rect 65566 25542 66424 25594
rect 63572 25520 66424 25542
rect 63954 25304 63960 25356
rect 64012 25344 64018 25356
rect 64325 25347 64383 25353
rect 64325 25344 64337 25347
rect 64012 25316 64337 25344
rect 64012 25304 64018 25316
rect 64325 25313 64337 25316
rect 64371 25313 64383 25347
rect 64325 25307 64383 25313
rect 64969 25347 65027 25353
rect 64969 25313 64981 25347
rect 65015 25344 65027 25347
rect 65429 25347 65487 25353
rect 65429 25344 65441 25347
rect 65015 25316 65441 25344
rect 65015 25313 65027 25316
rect 64969 25307 65027 25313
rect 65429 25313 65441 25316
rect 65475 25313 65487 25347
rect 65429 25307 65487 25313
rect 65058 25236 65064 25288
rect 65116 25236 65122 25288
rect 65150 25236 65156 25288
rect 65208 25236 65214 25288
rect 65794 25236 65800 25288
rect 65852 25276 65858 25288
rect 65981 25279 66039 25285
rect 65981 25276 65993 25279
rect 65852 25248 65993 25276
rect 65852 25236 65858 25248
rect 65981 25245 65993 25248
rect 66027 25245 66039 25279
rect 65981 25239 66039 25245
rect 64230 25100 64236 25152
rect 64288 25140 64294 25152
rect 64601 25143 64659 25149
rect 64601 25140 64613 25143
rect 64288 25112 64613 25140
rect 64288 25100 64294 25112
rect 64601 25109 64613 25112
rect 64647 25109 64659 25143
rect 64601 25103 64659 25109
rect 63572 25050 66424 25072
rect 63572 24998 64338 25050
rect 64390 24998 64402 25050
rect 64454 24998 64466 25050
rect 64518 24998 64530 25050
rect 64582 24998 64594 25050
rect 64646 24998 66424 25050
rect 63572 24976 66424 24998
rect 63865 24735 63923 24741
rect 63865 24701 63877 24735
rect 63911 24732 63923 24735
rect 64874 24732 64880 24744
rect 63911 24704 64880 24732
rect 63911 24701 63923 24704
rect 63865 24695 63923 24701
rect 64874 24692 64880 24704
rect 64932 24692 64938 24744
rect 63954 24556 63960 24608
rect 64012 24596 64018 24608
rect 65153 24599 65211 24605
rect 65153 24596 65165 24599
rect 64012 24568 65165 24596
rect 64012 24556 64018 24568
rect 65153 24565 65165 24568
rect 65199 24565 65211 24599
rect 65153 24559 65211 24565
rect 63572 24506 66424 24528
rect 63572 24454 65258 24506
rect 65310 24454 65322 24506
rect 65374 24454 65386 24506
rect 65438 24454 65450 24506
rect 65502 24454 65514 24506
rect 65566 24454 66424 24506
rect 63572 24432 66424 24454
rect 64230 24284 64236 24336
rect 64288 24324 64294 24336
rect 64325 24327 64383 24333
rect 64325 24324 64337 24327
rect 64288 24296 64337 24324
rect 64288 24284 64294 24296
rect 64325 24293 64337 24296
rect 64371 24293 64383 24327
rect 64325 24287 64383 24293
rect 64966 24284 64972 24336
rect 65024 24284 65030 24336
rect 63954 24148 63960 24200
rect 64012 24188 64018 24200
rect 64049 24191 64107 24197
rect 64049 24188 64061 24191
rect 64012 24160 64061 24188
rect 64012 24148 64018 24160
rect 64049 24157 64061 24160
rect 64095 24157 64107 24191
rect 64049 24151 64107 24157
rect 65794 24012 65800 24064
rect 65852 24012 65858 24064
rect 63572 23962 66424 23984
rect 63572 23910 64338 23962
rect 64390 23910 64402 23962
rect 64454 23910 64466 23962
rect 64518 23910 64530 23962
rect 64582 23910 64594 23962
rect 64646 23910 66424 23962
rect 63572 23888 66424 23910
rect 63034 23740 63040 23792
rect 63092 23780 63098 23792
rect 63862 23780 63868 23792
rect 63092 23752 63868 23780
rect 63092 23740 63098 23752
rect 63862 23740 63868 23752
rect 63920 23740 63926 23792
rect 62758 23604 62764 23656
rect 62816 23644 62822 23656
rect 63865 23647 63923 23653
rect 63865 23644 63877 23647
rect 62816 23616 63877 23644
rect 62816 23604 62822 23616
rect 63865 23613 63877 23616
rect 63911 23613 63923 23647
rect 63865 23607 63923 23613
rect 63402 23468 63408 23520
rect 63460 23508 63466 23520
rect 63678 23508 63684 23520
rect 63460 23480 63684 23508
rect 63460 23468 63466 23480
rect 63678 23468 63684 23480
rect 63736 23468 63742 23520
rect 64046 23468 64052 23520
rect 64104 23508 64110 23520
rect 65153 23511 65211 23517
rect 65153 23508 65165 23511
rect 64104 23480 65165 23508
rect 64104 23468 64110 23480
rect 65153 23477 65165 23480
rect 65199 23477 65211 23511
rect 65153 23471 65211 23477
rect 63572 23418 66424 23440
rect 63572 23366 65258 23418
rect 65310 23366 65322 23418
rect 65374 23366 65386 23418
rect 65438 23366 65450 23418
rect 65502 23366 65514 23418
rect 65566 23366 66424 23418
rect 63572 23344 66424 23366
rect 65058 23264 65064 23316
rect 65116 23304 65122 23316
rect 65245 23307 65303 23313
rect 65245 23304 65257 23307
rect 65116 23276 65257 23304
rect 65116 23264 65122 23276
rect 65245 23273 65257 23276
rect 65291 23273 65303 23307
rect 65245 23267 65303 23273
rect 64785 23239 64843 23245
rect 64785 23205 64797 23239
rect 64831 23236 64843 23239
rect 65978 23236 65984 23248
rect 64831 23208 65984 23236
rect 64831 23205 64843 23208
rect 64785 23199 64843 23205
rect 65978 23196 65984 23208
rect 66036 23196 66042 23248
rect 64046 23128 64052 23180
rect 64104 23128 64110 23180
rect 64877 23171 64935 23177
rect 64877 23137 64889 23171
rect 64923 23168 64935 23171
rect 64966 23168 64972 23180
rect 64923 23140 64972 23168
rect 64923 23137 64935 23140
rect 64877 23131 64935 23137
rect 64966 23128 64972 23140
rect 65024 23168 65030 23180
rect 66530 23168 66536 23180
rect 65024 23140 66536 23168
rect 65024 23128 65030 23140
rect 66530 23128 66536 23140
rect 66588 23128 66594 23180
rect 64693 23103 64751 23109
rect 64693 23069 64705 23103
rect 64739 23100 64751 23103
rect 65610 23100 65616 23112
rect 64739 23072 65616 23100
rect 64739 23069 64751 23072
rect 64693 23063 64751 23069
rect 65610 23060 65616 23072
rect 65668 23060 65674 23112
rect 63126 22992 63132 23044
rect 63184 23032 63190 23044
rect 64874 23032 64880 23044
rect 63184 23004 64880 23032
rect 63184 22992 63190 23004
rect 64874 22992 64880 23004
rect 64932 22992 64938 23044
rect 63572 22874 66424 22896
rect 63572 22822 64338 22874
rect 64390 22822 64402 22874
rect 64454 22822 64466 22874
rect 64518 22822 64530 22874
rect 64582 22822 64594 22874
rect 64646 22822 66424 22874
rect 63572 22800 66424 22822
rect 64601 22763 64659 22769
rect 64601 22729 64613 22763
rect 64647 22760 64659 22763
rect 64966 22760 64972 22772
rect 64647 22732 64972 22760
rect 64647 22729 64659 22732
rect 64601 22723 64659 22729
rect 64966 22720 64972 22732
rect 65024 22720 65030 22772
rect 63572 22330 66424 22352
rect 63572 22278 65258 22330
rect 65310 22278 65322 22330
rect 65374 22278 65386 22330
rect 65438 22278 65450 22330
rect 65502 22278 65514 22330
rect 65566 22278 66424 22330
rect 63572 22256 66424 22278
rect 65797 22219 65855 22225
rect 65797 22185 65809 22219
rect 65843 22216 65855 22219
rect 66346 22216 66352 22228
rect 65843 22188 66352 22216
rect 65843 22185 65855 22188
rect 65797 22179 65855 22185
rect 66346 22176 66352 22188
rect 66404 22176 66410 22228
rect 66162 22148 66168 22160
rect 65550 22120 66168 22148
rect 66162 22108 66168 22120
rect 66220 22108 66226 22160
rect 63954 21972 63960 22024
rect 64012 22012 64018 22024
rect 64049 22015 64107 22021
rect 64049 22012 64061 22015
rect 64012 21984 64061 22012
rect 64012 21972 64018 21984
rect 64049 21981 64061 21984
rect 64095 21981 64107 22015
rect 64049 21975 64107 21981
rect 64325 22015 64383 22021
rect 64325 21981 64337 22015
rect 64371 22012 64383 22015
rect 64690 22012 64696 22024
rect 64371 21984 64696 22012
rect 64371 21981 64383 21984
rect 64325 21975 64383 21981
rect 64690 21972 64696 21984
rect 64748 21972 64754 22024
rect 63572 21786 66424 21808
rect 63572 21734 64338 21786
rect 64390 21734 64402 21786
rect 64454 21734 64466 21786
rect 64518 21734 64530 21786
rect 64582 21734 64594 21786
rect 64646 21734 66424 21786
rect 63572 21712 66424 21734
rect 66073 21539 66131 21545
rect 66073 21505 66085 21539
rect 66119 21536 66131 21539
rect 66346 21536 66352 21548
rect 66119 21508 66352 21536
rect 66119 21505 66131 21508
rect 66073 21499 66131 21505
rect 66346 21496 66352 21508
rect 66404 21496 66410 21548
rect 63310 21428 63316 21480
rect 63368 21468 63374 21480
rect 63862 21468 63868 21480
rect 63368 21440 63868 21468
rect 63368 21428 63374 21440
rect 63862 21428 63868 21440
rect 63920 21468 63926 21480
rect 65061 21471 65119 21477
rect 65061 21468 65073 21471
rect 63920 21440 65073 21468
rect 63920 21428 63926 21440
rect 65061 21437 65073 21440
rect 65107 21437 65119 21471
rect 65061 21431 65119 21437
rect 65610 21400 65616 21412
rect 64892 21372 65616 21400
rect 64785 21335 64843 21341
rect 64785 21301 64797 21335
rect 64831 21332 64843 21335
rect 64892 21332 64920 21372
rect 65610 21360 65616 21372
rect 65668 21360 65674 21412
rect 64831 21304 64920 21332
rect 64831 21301 64843 21304
rect 64785 21295 64843 21301
rect 64966 21292 64972 21344
rect 65024 21332 65030 21344
rect 65429 21335 65487 21341
rect 65429 21332 65441 21335
rect 65024 21304 65441 21332
rect 65024 21292 65030 21304
rect 65429 21301 65441 21304
rect 65475 21301 65487 21335
rect 65429 21295 65487 21301
rect 63572 21242 66424 21264
rect 63572 21190 65258 21242
rect 65310 21190 65322 21242
rect 65374 21190 65386 21242
rect 65438 21190 65450 21242
rect 65502 21190 65514 21242
rect 65566 21190 66424 21242
rect 63572 21168 66424 21190
rect 64601 21131 64659 21137
rect 64601 21097 64613 21131
rect 64647 21128 64659 21131
rect 64690 21128 64696 21140
rect 64647 21100 64696 21128
rect 64647 21097 64659 21100
rect 64601 21091 64659 21097
rect 64690 21088 64696 21100
rect 64748 21088 64754 21140
rect 64966 21088 64972 21140
rect 65024 21088 65030 21140
rect 65061 21063 65119 21069
rect 65061 21029 65073 21063
rect 65107 21060 65119 21063
rect 65150 21060 65156 21072
rect 65107 21032 65156 21060
rect 65107 21029 65119 21032
rect 65061 21023 65119 21029
rect 65150 21020 65156 21032
rect 65208 21020 65214 21072
rect 65521 21063 65579 21069
rect 65521 21029 65533 21063
rect 65567 21060 65579 21063
rect 66070 21060 66076 21072
rect 65567 21032 66076 21060
rect 65567 21029 65579 21032
rect 65521 21023 65579 21029
rect 66070 21020 66076 21032
rect 66128 21020 66134 21072
rect 65245 20927 65303 20933
rect 65245 20893 65257 20927
rect 65291 20924 65303 20927
rect 65610 20924 65616 20936
rect 65291 20896 65616 20924
rect 65291 20893 65303 20896
rect 65245 20887 65303 20893
rect 65610 20884 65616 20896
rect 65668 20884 65674 20936
rect 65797 20791 65855 20797
rect 65797 20757 65809 20791
rect 65843 20788 65855 20791
rect 66162 20788 66168 20800
rect 65843 20760 66168 20788
rect 65843 20757 65855 20760
rect 65797 20751 65855 20757
rect 66162 20748 66168 20760
rect 66220 20748 66226 20800
rect 63572 20698 66424 20720
rect 63572 20646 64338 20698
rect 64390 20646 64402 20698
rect 64454 20646 64466 20698
rect 64518 20646 64530 20698
rect 64582 20646 64594 20698
rect 64646 20646 66424 20698
rect 63572 20624 66424 20646
rect 64138 20544 64144 20596
rect 64196 20584 64202 20596
rect 65886 20584 65892 20596
rect 64196 20556 65892 20584
rect 64196 20544 64202 20556
rect 65886 20544 65892 20556
rect 65944 20544 65950 20596
rect 64601 20519 64659 20525
rect 64601 20485 64613 20519
rect 64647 20516 64659 20519
rect 65058 20516 65064 20528
rect 64647 20488 65064 20516
rect 64647 20485 64659 20488
rect 64601 20479 64659 20485
rect 65058 20476 65064 20488
rect 65116 20476 65122 20528
rect 65245 20451 65303 20457
rect 65245 20417 65257 20451
rect 65291 20448 65303 20451
rect 65702 20448 65708 20460
rect 65291 20420 65708 20448
rect 65291 20417 65303 20420
rect 65245 20411 65303 20417
rect 65702 20408 65708 20420
rect 65760 20408 65766 20460
rect 65061 20383 65119 20389
rect 65061 20349 65073 20383
rect 65107 20380 65119 20383
rect 65794 20380 65800 20392
rect 65107 20352 65800 20380
rect 65107 20349 65119 20352
rect 65061 20343 65119 20349
rect 65794 20340 65800 20352
rect 65852 20340 65858 20392
rect 64966 20204 64972 20256
rect 65024 20204 65030 20256
rect 63572 20154 66424 20176
rect 63572 20102 65258 20154
rect 65310 20102 65322 20154
rect 65374 20102 65386 20154
rect 65438 20102 65450 20154
rect 65502 20102 65514 20154
rect 65566 20102 66424 20154
rect 63572 20080 66424 20102
rect 66162 19972 66168 19984
rect 65550 19944 66168 19972
rect 66162 19932 66168 19944
rect 66220 19932 66226 19984
rect 64046 19864 64052 19916
rect 64104 19864 64110 19916
rect 64325 19839 64383 19845
rect 64325 19805 64337 19839
rect 64371 19836 64383 19839
rect 64690 19836 64696 19848
rect 64371 19808 64696 19836
rect 64371 19805 64383 19808
rect 64325 19799 64383 19805
rect 64690 19796 64696 19808
rect 64748 19796 64754 19848
rect 65797 19703 65855 19709
rect 65797 19669 65809 19703
rect 65843 19700 65855 19703
rect 65978 19700 65984 19712
rect 65843 19672 65984 19700
rect 65843 19669 65855 19672
rect 65797 19663 65855 19669
rect 65978 19660 65984 19672
rect 66036 19660 66042 19712
rect 63572 19610 66424 19632
rect 63572 19558 64338 19610
rect 64390 19558 64402 19610
rect 64454 19558 64466 19610
rect 64518 19558 64530 19610
rect 64582 19558 64594 19610
rect 64646 19558 66424 19610
rect 63572 19536 66424 19558
rect 64601 19499 64659 19505
rect 64601 19465 64613 19499
rect 64647 19496 64659 19499
rect 64690 19496 64696 19508
rect 64647 19468 64696 19496
rect 64647 19465 64659 19468
rect 64601 19459 64659 19465
rect 64690 19456 64696 19468
rect 64748 19456 64754 19508
rect 65245 19363 65303 19369
rect 65245 19329 65257 19363
rect 65291 19360 65303 19363
rect 65610 19360 65616 19372
rect 65291 19332 65616 19360
rect 65291 19329 65303 19332
rect 65245 19323 65303 19329
rect 65610 19320 65616 19332
rect 65668 19320 65674 19372
rect 65058 19252 65064 19304
rect 65116 19252 65122 19304
rect 65978 19252 65984 19304
rect 66036 19252 66042 19304
rect 64969 19227 65027 19233
rect 64969 19193 64981 19227
rect 65015 19224 65027 19227
rect 65429 19227 65487 19233
rect 65429 19224 65441 19227
rect 65015 19196 65441 19224
rect 65015 19193 65027 19196
rect 64969 19187 65027 19193
rect 65429 19193 65441 19196
rect 65475 19193 65487 19227
rect 65429 19187 65487 19193
rect 63572 19066 66424 19088
rect 63572 19014 65258 19066
rect 65310 19014 65322 19066
rect 65374 19014 65386 19066
rect 65438 19014 65450 19066
rect 65502 19014 65514 19066
rect 65566 19014 66424 19066
rect 63572 18992 66424 19014
rect 64969 18819 65027 18825
rect 64969 18785 64981 18819
rect 65015 18816 65027 18819
rect 65429 18819 65487 18825
rect 65429 18816 65441 18819
rect 65015 18788 65441 18816
rect 65015 18785 65027 18788
rect 64969 18779 65027 18785
rect 65429 18785 65441 18788
rect 65475 18785 65487 18819
rect 65429 18779 65487 18785
rect 65058 18708 65064 18760
rect 65116 18708 65122 18760
rect 65245 18751 65303 18757
rect 65245 18717 65257 18751
rect 65291 18748 65303 18751
rect 65610 18748 65616 18760
rect 65291 18720 65616 18748
rect 65291 18717 65303 18720
rect 65245 18711 65303 18717
rect 65610 18708 65616 18720
rect 65668 18708 65674 18760
rect 65794 18708 65800 18760
rect 65852 18748 65858 18760
rect 65981 18751 66039 18757
rect 65981 18748 65993 18751
rect 65852 18720 65993 18748
rect 65852 18708 65858 18720
rect 65981 18717 65993 18720
rect 66027 18717 66039 18751
rect 65981 18711 66039 18717
rect 64601 18615 64659 18621
rect 64601 18581 64613 18615
rect 64647 18612 64659 18615
rect 64690 18612 64696 18624
rect 64647 18584 64696 18612
rect 64647 18581 64659 18584
rect 64601 18575 64659 18581
rect 64690 18572 64696 18584
rect 64748 18572 64754 18624
rect 63572 18522 66424 18544
rect 63572 18470 64338 18522
rect 64390 18470 64402 18522
rect 64454 18470 64466 18522
rect 64518 18470 64530 18522
rect 64582 18470 64594 18522
rect 64646 18470 66424 18522
rect 63572 18448 66424 18470
rect 64046 18232 64052 18284
rect 64104 18232 64110 18284
rect 64325 18275 64383 18281
rect 64325 18241 64337 18275
rect 64371 18272 64383 18275
rect 64690 18272 64696 18284
rect 64371 18244 64696 18272
rect 64371 18241 64383 18244
rect 64325 18235 64383 18241
rect 64690 18232 64696 18244
rect 64748 18232 64754 18284
rect 66162 18136 66168 18148
rect 65550 18108 66168 18136
rect 66162 18096 66168 18108
rect 66220 18096 66226 18148
rect 65794 18028 65800 18080
rect 65852 18028 65858 18080
rect 63572 17978 66424 18000
rect 63572 17926 65258 17978
rect 65310 17926 65322 17978
rect 65374 17926 65386 17978
rect 65438 17926 65450 17978
rect 65502 17926 65514 17978
rect 65566 17926 66424 17978
rect 63572 17904 66424 17926
rect 64230 17824 64236 17876
rect 64288 17864 64294 17876
rect 64877 17867 64935 17873
rect 64877 17864 64889 17867
rect 64288 17836 64889 17864
rect 64288 17824 64294 17836
rect 64877 17833 64889 17836
rect 64923 17833 64935 17867
rect 64877 17827 64935 17833
rect 65058 17824 65064 17876
rect 65116 17864 65122 17876
rect 65337 17867 65395 17873
rect 65337 17864 65349 17867
rect 65116 17836 65349 17864
rect 65116 17824 65122 17836
rect 65337 17833 65349 17836
rect 65383 17833 65395 17867
rect 65337 17827 65395 17833
rect 65705 17867 65763 17873
rect 65705 17833 65717 17867
rect 65751 17864 65763 17867
rect 66346 17864 66352 17876
rect 65751 17836 66352 17864
rect 65751 17833 65763 17836
rect 65705 17827 65763 17833
rect 66346 17824 66352 17836
rect 66404 17824 66410 17876
rect 64785 17799 64843 17805
rect 64785 17765 64797 17799
rect 64831 17796 64843 17799
rect 65794 17796 65800 17808
rect 64831 17768 65800 17796
rect 64831 17765 64843 17768
rect 64785 17759 64843 17765
rect 65794 17756 65800 17768
rect 65852 17756 65858 17808
rect 65702 17728 65708 17740
rect 64846 17700 65708 17728
rect 64846 17672 64874 17700
rect 65702 17688 65708 17700
rect 65760 17728 65766 17740
rect 65760 17700 65932 17728
rect 65760 17688 65766 17700
rect 64693 17663 64751 17669
rect 64693 17629 64705 17663
rect 64739 17660 64751 17663
rect 64846 17660 64880 17672
rect 64739 17632 64880 17660
rect 64739 17629 64751 17632
rect 64693 17623 64751 17629
rect 64874 17620 64880 17632
rect 64932 17620 64938 17672
rect 65904 17669 65932 17700
rect 65797 17663 65855 17669
rect 65797 17660 65809 17663
rect 65720 17632 65809 17660
rect 65720 17604 65748 17632
rect 65797 17629 65809 17632
rect 65843 17629 65855 17663
rect 65797 17623 65855 17629
rect 65889 17663 65947 17669
rect 65889 17629 65901 17663
rect 65935 17629 65947 17663
rect 65889 17623 65947 17629
rect 65150 17552 65156 17604
rect 65208 17592 65214 17604
rect 65245 17595 65303 17601
rect 65245 17592 65257 17595
rect 65208 17564 65257 17592
rect 65208 17552 65214 17564
rect 65245 17561 65257 17564
rect 65291 17561 65303 17595
rect 65245 17555 65303 17561
rect 65702 17552 65708 17604
rect 65760 17552 65766 17604
rect 63572 17434 66424 17456
rect 63572 17382 64338 17434
rect 64390 17382 64402 17434
rect 64454 17382 64466 17434
rect 64518 17382 64530 17434
rect 64582 17382 64594 17434
rect 64646 17382 66424 17434
rect 63572 17360 66424 17382
rect 64230 17280 64236 17332
rect 64288 17320 64294 17332
rect 64509 17323 64567 17329
rect 64509 17320 64521 17323
rect 64288 17292 64521 17320
rect 64288 17280 64294 17292
rect 64509 17289 64521 17292
rect 64555 17289 64567 17323
rect 64509 17283 64567 17289
rect 63572 16890 66424 16912
rect 63572 16838 65258 16890
rect 65310 16838 65322 16890
rect 65374 16838 65386 16890
rect 65438 16838 65450 16890
rect 65502 16838 65514 16890
rect 65566 16838 66424 16890
rect 63572 16816 66424 16838
rect 64966 16736 64972 16788
rect 65024 16736 65030 16788
rect 64984 16708 65012 16736
rect 65150 16708 65156 16720
rect 64984 16680 65156 16708
rect 64984 16640 65012 16680
rect 65150 16668 65156 16680
rect 65208 16668 65214 16720
rect 65429 16643 65487 16649
rect 65429 16640 65441 16643
rect 64984 16612 65441 16640
rect 65429 16609 65441 16612
rect 65475 16609 65487 16643
rect 65429 16603 65487 16609
rect 63310 16396 63316 16448
rect 63368 16436 63374 16448
rect 65886 16436 65892 16448
rect 63368 16408 65892 16436
rect 63368 16396 63374 16408
rect 65886 16396 65892 16408
rect 65944 16396 65950 16448
rect 66070 16396 66076 16448
rect 66128 16396 66134 16448
rect 63572 16346 66424 16368
rect 63572 16294 64338 16346
rect 64390 16294 64402 16346
rect 64454 16294 64466 16346
rect 64518 16294 64530 16346
rect 64582 16294 64594 16346
rect 64646 16294 66424 16346
rect 63572 16272 66424 16294
rect 64874 16232 64880 16244
rect 64708 16204 64880 16232
rect 64708 16105 64736 16204
rect 64874 16192 64880 16204
rect 64932 16192 64938 16244
rect 64782 16124 64788 16176
rect 64840 16164 64846 16176
rect 65337 16167 65395 16173
rect 65337 16164 65349 16167
rect 64840 16136 65349 16164
rect 64840 16124 64846 16136
rect 65337 16133 65349 16136
rect 65383 16133 65395 16167
rect 65978 16164 65984 16176
rect 65337 16127 65395 16133
rect 65444 16136 65984 16164
rect 64693 16099 64751 16105
rect 64693 16065 64705 16099
rect 64739 16065 64751 16099
rect 64693 16059 64751 16065
rect 64598 15988 64604 16040
rect 64656 16028 64662 16040
rect 64877 16031 64935 16037
rect 64877 16028 64889 16031
rect 64656 16000 64889 16028
rect 64656 15988 64662 16000
rect 64877 15997 64889 16000
rect 64923 15997 64935 16031
rect 65444 16028 65472 16136
rect 65978 16124 65984 16136
rect 66036 16124 66042 16176
rect 65886 16056 65892 16108
rect 65944 16096 65950 16108
rect 66438 16096 66444 16108
rect 65944 16068 66444 16096
rect 65944 16056 65950 16068
rect 66438 16056 66444 16068
rect 66496 16056 66502 16108
rect 64877 15991 64935 15997
rect 65168 16000 65472 16028
rect 65705 16031 65763 16037
rect 64785 15895 64843 15901
rect 64785 15861 64797 15895
rect 64831 15892 64843 15895
rect 65168 15892 65196 16000
rect 65705 15997 65717 16031
rect 65751 16028 65763 16031
rect 66070 16028 66076 16040
rect 65751 16000 66076 16028
rect 65751 15997 65763 16000
rect 65705 15991 65763 15997
rect 66070 15988 66076 16000
rect 66128 15988 66134 16040
rect 65797 15963 65855 15969
rect 65797 15960 65809 15963
rect 65260 15932 65809 15960
rect 65260 15901 65288 15932
rect 65797 15929 65809 15932
rect 65843 15929 65855 15963
rect 65797 15923 65855 15929
rect 64831 15864 65196 15892
rect 65245 15895 65303 15901
rect 64831 15861 64843 15864
rect 64785 15855 64843 15861
rect 65245 15861 65257 15895
rect 65291 15861 65303 15895
rect 65245 15855 65303 15861
rect 63572 15802 66424 15824
rect 63572 15750 65258 15802
rect 65310 15750 65322 15802
rect 65374 15750 65386 15802
rect 65438 15750 65450 15802
rect 65502 15750 65514 15802
rect 65566 15750 66424 15802
rect 63572 15728 66424 15750
rect 64598 15648 64604 15700
rect 64656 15648 64662 15700
rect 62758 15308 62764 15360
rect 62816 15348 62822 15360
rect 64138 15348 64144 15360
rect 62816 15320 64144 15348
rect 62816 15308 62822 15320
rect 64138 15308 64144 15320
rect 64196 15308 64202 15360
rect 63572 15258 66424 15280
rect 63572 15206 64338 15258
rect 64390 15206 64402 15258
rect 64454 15206 64466 15258
rect 64518 15206 64530 15258
rect 64582 15206 64594 15258
rect 64646 15206 66424 15258
rect 63572 15184 66424 15206
rect 64325 15011 64383 15017
rect 64325 14977 64337 15011
rect 64371 15008 64383 15011
rect 64782 15008 64788 15020
rect 64371 14980 64788 15008
rect 64371 14977 64383 14980
rect 64325 14971 64383 14977
rect 64782 14968 64788 14980
rect 64840 14968 64846 15020
rect 63862 14900 63868 14952
rect 63920 14940 63926 14952
rect 64049 14943 64107 14949
rect 64049 14940 64061 14943
rect 63920 14912 64061 14940
rect 63920 14900 63926 14912
rect 64049 14909 64061 14912
rect 64095 14909 64107 14943
rect 64049 14903 64107 14909
rect 65058 14832 65064 14884
rect 65116 14832 65122 14884
rect 62942 14764 62948 14816
rect 63000 14804 63006 14816
rect 63678 14804 63684 14816
rect 63000 14776 63684 14804
rect 63000 14764 63006 14776
rect 63678 14764 63684 14776
rect 63736 14764 63742 14816
rect 65150 14764 65156 14816
rect 65208 14804 65214 14816
rect 65794 14804 65800 14816
rect 65208 14776 65800 14804
rect 65208 14764 65214 14776
rect 65794 14764 65800 14776
rect 65852 14764 65858 14816
rect 63572 14714 66424 14736
rect 63572 14662 65258 14714
rect 65310 14662 65322 14714
rect 65374 14662 65386 14714
rect 65438 14662 65450 14714
rect 65502 14662 65514 14714
rect 65566 14662 66424 14714
rect 63572 14640 66424 14662
rect 63572 14170 66424 14192
rect 63572 14118 64338 14170
rect 64390 14118 64402 14170
rect 64454 14118 64466 14170
rect 64518 14118 64530 14170
rect 64582 14118 64594 14170
rect 64646 14118 66424 14170
rect 63572 14096 66424 14118
rect 63034 13812 63040 13864
rect 63092 13852 63098 13864
rect 63586 13852 63592 13864
rect 63092 13824 63592 13852
rect 63092 13812 63098 13824
rect 63586 13812 63592 13824
rect 63644 13812 63650 13864
rect 63572 13626 66424 13648
rect 63572 13574 65258 13626
rect 65310 13574 65322 13626
rect 65374 13574 65386 13626
rect 65438 13574 65450 13626
rect 65502 13574 65514 13626
rect 65566 13574 66424 13626
rect 63572 13552 66424 13574
rect 65702 13472 65708 13524
rect 65760 13512 65766 13524
rect 65797 13515 65855 13521
rect 65797 13512 65809 13515
rect 65760 13484 65809 13512
rect 65760 13472 65766 13484
rect 65797 13481 65809 13484
rect 65843 13481 65855 13515
rect 65797 13475 65855 13481
rect 64230 13404 64236 13456
rect 64288 13444 64294 13456
rect 64325 13447 64383 13453
rect 64325 13444 64337 13447
rect 64288 13416 64337 13444
rect 64288 13404 64294 13416
rect 64325 13413 64337 13416
rect 64371 13413 64383 13447
rect 65610 13444 65616 13456
rect 65550 13416 65616 13444
rect 64325 13407 64383 13413
rect 65610 13404 65616 13416
rect 65668 13444 65674 13456
rect 66162 13444 66168 13456
rect 65668 13416 66168 13444
rect 65668 13404 65674 13416
rect 66162 13404 66168 13416
rect 66220 13404 66226 13456
rect 63862 13268 63868 13320
rect 63920 13308 63926 13320
rect 64049 13311 64107 13317
rect 64049 13308 64061 13311
rect 63920 13280 64061 13308
rect 63920 13268 63926 13280
rect 64049 13277 64061 13280
rect 64095 13277 64107 13311
rect 64049 13271 64107 13277
rect 63572 13082 66424 13104
rect 63572 13030 64338 13082
rect 64390 13030 64402 13082
rect 64454 13030 64466 13082
rect 64518 13030 64530 13082
rect 64582 13030 64594 13082
rect 64646 13030 66424 13082
rect 63572 13008 66424 13030
rect 65702 12792 65708 12844
rect 65760 12832 65766 12844
rect 65981 12835 66039 12841
rect 65981 12832 65993 12835
rect 65760 12804 65993 12832
rect 65760 12792 65766 12804
rect 65981 12801 65993 12804
rect 66027 12801 66039 12835
rect 65981 12795 66039 12801
rect 64966 12588 64972 12640
rect 65024 12628 65030 12640
rect 65429 12631 65487 12637
rect 65429 12628 65441 12631
rect 65024 12600 65441 12628
rect 65024 12588 65030 12600
rect 65429 12597 65441 12600
rect 65475 12597 65487 12631
rect 65429 12591 65487 12597
rect 63572 12538 66424 12560
rect 63572 12486 65258 12538
rect 65310 12486 65322 12538
rect 65374 12486 65386 12538
rect 65438 12486 65450 12538
rect 65502 12486 65514 12538
rect 65566 12486 66424 12538
rect 63572 12464 66424 12486
rect 65610 12356 65616 12368
rect 65550 12328 65616 12356
rect 65610 12316 65616 12328
rect 65668 12316 65674 12368
rect 63862 12180 63868 12232
rect 63920 12220 63926 12232
rect 64049 12223 64107 12229
rect 64049 12220 64061 12223
rect 63920 12192 64061 12220
rect 63920 12180 63926 12192
rect 64049 12189 64061 12192
rect 64095 12189 64107 12223
rect 64049 12183 64107 12189
rect 64325 12223 64383 12229
rect 64325 12189 64337 12223
rect 64371 12220 64383 12223
rect 64690 12220 64696 12232
rect 64371 12192 64696 12220
rect 64371 12189 64383 12192
rect 64325 12183 64383 12189
rect 64690 12180 64696 12192
rect 64748 12180 64754 12232
rect 66073 12223 66131 12229
rect 66073 12189 66085 12223
rect 66119 12220 66131 12223
rect 66346 12220 66352 12232
rect 66119 12192 66352 12220
rect 66119 12189 66131 12192
rect 66073 12183 66131 12189
rect 66346 12180 66352 12192
rect 66404 12180 66410 12232
rect 63572 11994 66424 12016
rect 63572 11942 64338 11994
rect 64390 11942 64402 11994
rect 64454 11942 64466 11994
rect 64518 11942 64530 11994
rect 64582 11942 64594 11994
rect 64646 11942 66424 11994
rect 63572 11920 66424 11942
rect 64230 11840 64236 11892
rect 64288 11880 64294 11892
rect 64601 11883 64659 11889
rect 64601 11880 64613 11883
rect 64288 11852 64613 11880
rect 64288 11840 64294 11852
rect 64601 11849 64613 11852
rect 64647 11849 64659 11883
rect 64601 11843 64659 11849
rect 65150 11704 65156 11756
rect 65208 11704 65214 11756
rect 64966 11636 64972 11688
rect 65024 11636 65030 11688
rect 63954 11500 63960 11552
rect 64012 11540 64018 11552
rect 65061 11543 65119 11549
rect 65061 11540 65073 11543
rect 64012 11512 65073 11540
rect 64012 11500 64018 11512
rect 65061 11509 65073 11512
rect 65107 11509 65119 11543
rect 65061 11503 65119 11509
rect 63572 11450 66424 11472
rect 63572 11398 65258 11450
rect 65310 11398 65322 11450
rect 65374 11398 65386 11450
rect 65438 11398 65450 11450
rect 65502 11398 65514 11450
rect 65566 11398 66424 11450
rect 63572 11376 66424 11398
rect 64509 11339 64567 11345
rect 64509 11305 64521 11339
rect 64555 11336 64567 11339
rect 64690 11336 64696 11348
rect 64555 11308 64696 11336
rect 64555 11305 64567 11308
rect 64509 11299 64567 11305
rect 64690 11296 64696 11308
rect 64748 11296 64754 11348
rect 63678 11228 63684 11280
rect 63736 11268 63742 11280
rect 64877 11271 64935 11277
rect 64877 11268 64889 11271
rect 63736 11240 64889 11268
rect 63736 11228 63742 11240
rect 64877 11237 64889 11240
rect 64923 11268 64935 11271
rect 66346 11268 66352 11280
rect 64923 11240 66352 11268
rect 64923 11237 64935 11240
rect 64877 11231 64935 11237
rect 66346 11228 66352 11240
rect 66404 11228 66410 11280
rect 64969 11203 65027 11209
rect 64969 11169 64981 11203
rect 65015 11200 65027 11203
rect 66162 11200 66168 11212
rect 65015 11172 66168 11200
rect 65015 11169 65027 11172
rect 64969 11163 65027 11169
rect 66162 11160 66168 11172
rect 66220 11160 66226 11212
rect 65150 11092 65156 11144
rect 65208 11092 65214 11144
rect 63572 10906 66424 10928
rect 63572 10854 64338 10906
rect 64390 10854 64402 10906
rect 64454 10854 64466 10906
rect 64518 10854 64530 10906
rect 64582 10854 64594 10906
rect 64646 10854 66424 10906
rect 63572 10832 66424 10854
rect 64874 10616 64880 10668
rect 64932 10656 64938 10668
rect 65153 10659 65211 10665
rect 65153 10656 65165 10659
rect 64932 10628 65165 10656
rect 64932 10616 64938 10628
rect 65153 10625 65165 10628
rect 65199 10625 65211 10659
rect 65153 10619 65211 10625
rect 65061 10591 65119 10597
rect 65061 10557 65073 10591
rect 65107 10588 65119 10591
rect 65794 10588 65800 10600
rect 65107 10560 65800 10588
rect 65107 10557 65119 10560
rect 65061 10551 65119 10557
rect 65794 10548 65800 10560
rect 65852 10548 65858 10600
rect 64601 10455 64659 10461
rect 64601 10421 64613 10455
rect 64647 10452 64659 10455
rect 64782 10452 64788 10464
rect 64647 10424 64788 10452
rect 64647 10421 64659 10424
rect 64601 10415 64659 10421
rect 64782 10412 64788 10424
rect 64840 10412 64846 10464
rect 64874 10412 64880 10464
rect 64932 10452 64938 10464
rect 64969 10455 65027 10461
rect 64969 10452 64981 10455
rect 64932 10424 64981 10452
rect 64932 10412 64938 10424
rect 64969 10421 64981 10424
rect 65015 10421 65027 10455
rect 64969 10415 65027 10421
rect 63572 10362 66424 10384
rect 63572 10310 65258 10362
rect 65310 10310 65322 10362
rect 65374 10310 65386 10362
rect 65438 10310 65450 10362
rect 65502 10310 65514 10362
rect 65566 10310 66424 10362
rect 63572 10288 66424 10310
rect 64969 10251 65027 10257
rect 64969 10217 64981 10251
rect 65015 10248 65027 10251
rect 65702 10248 65708 10260
rect 65015 10220 65708 10248
rect 65015 10217 65027 10220
rect 64969 10211 65027 10217
rect 65702 10208 65708 10220
rect 65760 10208 65766 10260
rect 64966 10112 64972 10124
rect 64800 10084 64972 10112
rect 64800 10053 64828 10084
rect 64966 10072 64972 10084
rect 65024 10072 65030 10124
rect 64785 10047 64843 10053
rect 64785 10013 64797 10047
rect 64831 10013 64843 10047
rect 64785 10007 64843 10013
rect 64874 10004 64880 10056
rect 64932 10044 64938 10056
rect 65978 10044 65984 10056
rect 64932 10016 65984 10044
rect 64932 10004 64938 10016
rect 65978 10004 65984 10016
rect 66036 10004 66042 10056
rect 65337 9911 65395 9917
rect 65337 9877 65349 9911
rect 65383 9908 65395 9911
rect 65702 9908 65708 9920
rect 65383 9880 65708 9908
rect 65383 9877 65395 9880
rect 65337 9871 65395 9877
rect 65702 9868 65708 9880
rect 65760 9868 65766 9920
rect 63572 9818 66424 9840
rect 63572 9766 64338 9818
rect 64390 9766 64402 9818
rect 64454 9766 64466 9818
rect 64518 9766 64530 9818
rect 64582 9766 64594 9818
rect 64646 9766 66424 9818
rect 63572 9744 66424 9766
rect 65794 9460 65800 9512
rect 65852 9500 65858 9512
rect 65981 9503 66039 9509
rect 65981 9500 65993 9503
rect 65852 9472 65993 9500
rect 65852 9460 65858 9472
rect 65981 9469 65993 9472
rect 66027 9469 66039 9503
rect 65981 9463 66039 9469
rect 64966 9324 64972 9376
rect 65024 9364 65030 9376
rect 65429 9367 65487 9373
rect 65429 9364 65441 9367
rect 65024 9336 65441 9364
rect 65024 9324 65030 9336
rect 65429 9333 65441 9336
rect 65475 9333 65487 9367
rect 65429 9327 65487 9333
rect 63572 9274 66424 9296
rect 63572 9222 65258 9274
rect 65310 9222 65322 9274
rect 65374 9222 65386 9274
rect 65438 9222 65450 9274
rect 65502 9222 65514 9274
rect 65566 9222 66424 9274
rect 63572 9200 66424 9222
rect 65610 9092 65616 9104
rect 65550 9064 65616 9092
rect 65610 9052 65616 9064
rect 65668 9052 65674 9104
rect 63862 8916 63868 8968
rect 63920 8956 63926 8968
rect 64049 8959 64107 8965
rect 64049 8956 64061 8959
rect 63920 8928 64061 8956
rect 63920 8916 63926 8928
rect 64049 8925 64061 8928
rect 64095 8925 64107 8959
rect 64049 8919 64107 8925
rect 64325 8959 64383 8965
rect 64325 8925 64337 8959
rect 64371 8956 64383 8959
rect 64690 8956 64696 8968
rect 64371 8928 64696 8956
rect 64371 8925 64383 8928
rect 64325 8919 64383 8925
rect 64690 8916 64696 8928
rect 64748 8916 64754 8968
rect 65797 8823 65855 8829
rect 65797 8789 65809 8823
rect 65843 8820 65855 8823
rect 65978 8820 65984 8832
rect 65843 8792 65984 8820
rect 65843 8789 65855 8792
rect 65797 8783 65855 8789
rect 65978 8780 65984 8792
rect 66036 8780 66042 8832
rect 63572 8730 66424 8752
rect 63572 8678 64338 8730
rect 64390 8678 64402 8730
rect 64454 8678 64466 8730
rect 64518 8678 64530 8730
rect 64582 8678 64594 8730
rect 64646 8678 66424 8730
rect 63572 8656 66424 8678
rect 64601 8619 64659 8625
rect 64601 8585 64613 8619
rect 64647 8616 64659 8619
rect 64690 8616 64696 8628
rect 64647 8588 64696 8616
rect 64647 8585 64659 8588
rect 64601 8579 64659 8585
rect 64690 8576 64696 8588
rect 64748 8576 64754 8628
rect 65242 8440 65248 8492
rect 65300 8480 65306 8492
rect 65886 8480 65892 8492
rect 65300 8452 65892 8480
rect 65300 8440 65306 8452
rect 65886 8440 65892 8452
rect 65944 8440 65950 8492
rect 65978 8440 65984 8492
rect 66036 8440 66042 8492
rect 65058 8372 65064 8424
rect 65116 8372 65122 8424
rect 64969 8347 65027 8353
rect 64969 8313 64981 8347
rect 65015 8344 65027 8347
rect 65429 8347 65487 8353
rect 65429 8344 65441 8347
rect 65015 8316 65441 8344
rect 65015 8313 65027 8316
rect 64969 8307 65027 8313
rect 65429 8313 65441 8316
rect 65475 8313 65487 8347
rect 65429 8307 65487 8313
rect 63572 8186 66424 8208
rect 63572 8134 65258 8186
rect 65310 8134 65322 8186
rect 65374 8134 65386 8186
rect 65438 8134 65450 8186
rect 65502 8134 65514 8186
rect 65566 8134 66424 8186
rect 63572 8112 66424 8134
rect 65794 8032 65800 8084
rect 65852 8032 65858 8084
rect 65610 8004 65616 8016
rect 65550 7976 65616 8004
rect 65610 7964 65616 7976
rect 65668 8004 65674 8016
rect 66070 8004 66076 8016
rect 65668 7976 66076 8004
rect 65668 7964 65674 7976
rect 66070 7964 66076 7976
rect 66128 7964 66134 8016
rect 64046 7896 64052 7948
rect 64104 7896 64110 7948
rect 64325 7871 64383 7877
rect 64325 7837 64337 7871
rect 64371 7868 64383 7871
rect 64690 7868 64696 7880
rect 64371 7840 64696 7868
rect 64371 7837 64383 7840
rect 64325 7831 64383 7837
rect 64690 7828 64696 7840
rect 64748 7828 64754 7880
rect 63572 7642 66424 7664
rect 63572 7590 64338 7642
rect 64390 7590 64402 7642
rect 64454 7590 64466 7642
rect 64518 7590 64530 7642
rect 64582 7590 64594 7642
rect 64646 7590 66424 7642
rect 63572 7568 66424 7590
rect 64138 7488 64144 7540
rect 64196 7528 64202 7540
rect 64417 7531 64475 7537
rect 64417 7528 64429 7531
rect 64196 7500 64429 7528
rect 64196 7488 64202 7500
rect 64417 7497 64429 7500
rect 64463 7497 64475 7531
rect 64417 7491 64475 7497
rect 64601 7531 64659 7537
rect 64601 7497 64613 7531
rect 64647 7528 64659 7531
rect 64690 7528 64696 7540
rect 64647 7500 64696 7528
rect 64647 7497 64659 7500
rect 64601 7491 64659 7497
rect 64690 7488 64696 7500
rect 64748 7488 64754 7540
rect 64782 7352 64788 7404
rect 64840 7392 64846 7404
rect 65061 7395 65119 7401
rect 65061 7392 65073 7395
rect 64840 7364 65073 7392
rect 64840 7352 64846 7364
rect 65061 7361 65073 7364
rect 65107 7361 65119 7395
rect 65061 7355 65119 7361
rect 65245 7395 65303 7401
rect 65245 7361 65257 7395
rect 65291 7392 65303 7395
rect 65886 7392 65892 7404
rect 65291 7364 65892 7392
rect 65291 7361 65303 7364
rect 65245 7355 65303 7361
rect 65886 7352 65892 7364
rect 65944 7352 65950 7404
rect 64966 7284 64972 7336
rect 65024 7284 65030 7336
rect 65978 7284 65984 7336
rect 66036 7284 66042 7336
rect 65429 7191 65487 7197
rect 65429 7157 65441 7191
rect 65475 7188 65487 7191
rect 65610 7188 65616 7200
rect 65475 7160 65616 7188
rect 65475 7157 65487 7160
rect 65429 7151 65487 7157
rect 65610 7148 65616 7160
rect 65668 7148 65674 7200
rect 63572 7098 66424 7120
rect 63572 7046 65258 7098
rect 65310 7046 65322 7098
rect 65374 7046 65386 7098
rect 65438 7046 65450 7098
rect 65502 7046 65514 7098
rect 65566 7046 66424 7098
rect 63572 7024 66424 7046
rect 64138 6944 64144 6996
rect 64196 6984 64202 6996
rect 64785 6987 64843 6993
rect 64785 6984 64797 6987
rect 64196 6956 64797 6984
rect 64196 6944 64202 6956
rect 64785 6953 64797 6956
rect 64831 6953 64843 6987
rect 64785 6947 64843 6953
rect 65610 6944 65616 6996
rect 65668 6944 65674 6996
rect 65794 6916 65800 6928
rect 65536 6888 65800 6916
rect 63770 6808 63776 6860
rect 63828 6848 63834 6860
rect 63865 6851 63923 6857
rect 63865 6848 63877 6851
rect 63828 6820 63877 6848
rect 63828 6808 63834 6820
rect 63865 6817 63877 6820
rect 63911 6817 63923 6851
rect 63865 6811 63923 6817
rect 64693 6851 64751 6857
rect 64693 6817 64705 6851
rect 64739 6848 64751 6851
rect 65536 6848 65564 6888
rect 65794 6876 65800 6888
rect 65852 6876 65858 6928
rect 64739 6820 65564 6848
rect 64739 6817 64751 6820
rect 64693 6811 64751 6817
rect 65702 6808 65708 6860
rect 65760 6808 65766 6860
rect 64141 6783 64199 6789
rect 64141 6749 64153 6783
rect 64187 6780 64199 6783
rect 64601 6783 64659 6789
rect 64601 6780 64613 6783
rect 64187 6752 64613 6780
rect 64187 6749 64199 6752
rect 64141 6743 64199 6749
rect 64601 6749 64613 6752
rect 64647 6780 64659 6783
rect 64874 6780 64880 6792
rect 64647 6752 64880 6780
rect 64647 6749 64659 6752
rect 64601 6743 64659 6749
rect 64874 6740 64880 6752
rect 64932 6740 64938 6792
rect 65794 6740 65800 6792
rect 65852 6740 65858 6792
rect 65058 6672 65064 6724
rect 65116 6712 65122 6724
rect 65153 6715 65211 6721
rect 65153 6712 65165 6715
rect 65116 6684 65165 6712
rect 65116 6672 65122 6684
rect 65153 6681 65165 6684
rect 65199 6681 65211 6715
rect 65153 6675 65211 6681
rect 64230 6604 64236 6656
rect 64288 6644 64294 6656
rect 65245 6647 65303 6653
rect 65245 6644 65257 6647
rect 64288 6616 65257 6644
rect 64288 6604 64294 6616
rect 65245 6613 65257 6616
rect 65291 6613 65303 6647
rect 65245 6607 65303 6613
rect 63572 6554 66424 6576
rect 63572 6502 64338 6554
rect 64390 6502 64402 6554
rect 64454 6502 64466 6554
rect 64518 6502 64530 6554
rect 64582 6502 64594 6554
rect 64646 6502 66424 6554
rect 63572 6480 66424 6502
rect 64138 6400 64144 6452
rect 64196 6440 64202 6452
rect 64417 6443 64475 6449
rect 64417 6440 64429 6443
rect 64196 6412 64429 6440
rect 64196 6400 64202 6412
rect 64417 6409 64429 6412
rect 64463 6409 64475 6443
rect 64417 6403 64475 6409
rect 63954 6332 63960 6384
rect 64012 6372 64018 6384
rect 64693 6375 64751 6381
rect 64693 6372 64705 6375
rect 64012 6344 64705 6372
rect 64012 6332 64018 6344
rect 64693 6341 64705 6344
rect 64739 6341 64751 6375
rect 64693 6335 64751 6341
rect 64874 6264 64880 6316
rect 64932 6304 64938 6316
rect 65245 6307 65303 6313
rect 65245 6304 65257 6307
rect 64932 6276 65257 6304
rect 64932 6264 64938 6276
rect 65245 6273 65257 6276
rect 65291 6273 65303 6307
rect 65245 6267 65303 6273
rect 65153 6239 65211 6245
rect 65153 6205 65165 6239
rect 65199 6236 65211 6239
rect 65978 6236 65984 6248
rect 65199 6208 65984 6236
rect 65199 6205 65211 6208
rect 65153 6199 65211 6205
rect 65978 6196 65984 6208
rect 66036 6196 66042 6248
rect 64690 6060 64696 6112
rect 64748 6100 64754 6112
rect 65061 6103 65119 6109
rect 65061 6100 65073 6103
rect 64748 6072 65073 6100
rect 64748 6060 64754 6072
rect 65061 6069 65073 6072
rect 65107 6069 65119 6103
rect 65061 6063 65119 6069
rect 63572 6010 66424 6032
rect 63572 5958 65258 6010
rect 65310 5958 65322 6010
rect 65374 5958 65386 6010
rect 65438 5958 65450 6010
rect 65502 5958 65514 6010
rect 65566 5958 66424 6010
rect 63572 5936 66424 5958
rect 64138 5856 64144 5908
rect 64196 5856 64202 5908
rect 64690 5856 64696 5908
rect 64748 5856 64754 5908
rect 64874 5856 64880 5908
rect 64932 5896 64938 5908
rect 65426 5896 65432 5908
rect 64932 5868 65432 5896
rect 64932 5856 64938 5868
rect 65426 5856 65432 5868
rect 65484 5896 65490 5908
rect 65794 5896 65800 5908
rect 65484 5868 65800 5896
rect 65484 5856 65490 5868
rect 65794 5856 65800 5868
rect 65852 5856 65858 5908
rect 64233 5831 64291 5837
rect 64233 5797 64245 5831
rect 64279 5828 64291 5831
rect 65702 5828 65708 5840
rect 64279 5800 65708 5828
rect 64279 5797 64291 5800
rect 64233 5791 64291 5797
rect 65702 5788 65708 5800
rect 65760 5788 65766 5840
rect 64782 5760 64788 5772
rect 64064 5732 64788 5760
rect 63954 5652 63960 5704
rect 64012 5692 64018 5704
rect 64064 5701 64092 5732
rect 64782 5720 64788 5732
rect 64840 5720 64846 5772
rect 65058 5720 65064 5772
rect 65116 5760 65122 5772
rect 65245 5763 65303 5769
rect 65245 5760 65257 5763
rect 65116 5732 65257 5760
rect 65116 5720 65122 5732
rect 65245 5729 65257 5732
rect 65291 5729 65303 5763
rect 65245 5723 65303 5729
rect 64049 5695 64107 5701
rect 64049 5692 64061 5695
rect 64012 5664 64061 5692
rect 64012 5652 64018 5664
rect 64049 5661 64061 5664
rect 64095 5661 64107 5695
rect 64049 5655 64107 5661
rect 64690 5652 64696 5704
rect 64748 5692 64754 5704
rect 65337 5695 65395 5701
rect 65337 5692 65349 5695
rect 64748 5664 65349 5692
rect 64748 5652 64754 5664
rect 65337 5661 65349 5664
rect 65383 5661 65395 5695
rect 65337 5655 65395 5661
rect 65426 5652 65432 5704
rect 65484 5652 65490 5704
rect 64601 5627 64659 5633
rect 64601 5593 64613 5627
rect 64647 5624 64659 5627
rect 64966 5624 64972 5636
rect 64647 5596 64972 5624
rect 64647 5593 64659 5596
rect 64601 5587 64659 5593
rect 64966 5584 64972 5596
rect 65024 5584 65030 5636
rect 64782 5516 64788 5568
rect 64840 5556 64846 5568
rect 64877 5559 64935 5565
rect 64877 5556 64889 5559
rect 64840 5528 64889 5556
rect 64840 5516 64846 5528
rect 64877 5525 64889 5528
rect 64923 5525 64935 5559
rect 64877 5519 64935 5525
rect 63572 5466 66424 5488
rect 63572 5414 64338 5466
rect 64390 5414 64402 5466
rect 64454 5414 64466 5466
rect 64518 5414 64530 5466
rect 64582 5414 64594 5466
rect 64646 5414 66424 5466
rect 63572 5392 66424 5414
rect 63862 5176 63868 5228
rect 63920 5176 63926 5228
rect 64141 5219 64199 5225
rect 64141 5185 64153 5219
rect 64187 5216 64199 5219
rect 64782 5216 64788 5228
rect 64187 5188 64788 5216
rect 64187 5185 64199 5188
rect 64141 5179 64199 5185
rect 64782 5176 64788 5188
rect 64840 5176 64846 5228
rect 65610 5148 65616 5160
rect 65274 5120 65616 5148
rect 65610 5108 65616 5120
rect 65668 5148 65674 5160
rect 66070 5148 66076 5160
rect 65668 5120 66076 5148
rect 65668 5108 65674 5120
rect 66070 5108 66076 5120
rect 66128 5108 66134 5160
rect 65613 5015 65671 5021
rect 65613 4981 65625 5015
rect 65659 5012 65671 5015
rect 65702 5012 65708 5024
rect 65659 4984 65708 5012
rect 65659 4981 65671 4984
rect 65613 4975 65671 4981
rect 65702 4972 65708 4984
rect 65760 4972 65766 5024
rect 63572 4922 66424 4944
rect 63572 4870 65258 4922
rect 65310 4870 65322 4922
rect 65374 4870 65386 4922
rect 65438 4870 65450 4922
rect 65502 4870 65514 4922
rect 65566 4870 66424 4922
rect 63572 4848 66424 4870
rect 65797 4811 65855 4817
rect 65797 4777 65809 4811
rect 65843 4808 65855 4811
rect 65978 4808 65984 4820
rect 65843 4780 65984 4808
rect 65843 4777 65855 4780
rect 65797 4771 65855 4777
rect 65978 4768 65984 4780
rect 66036 4768 66042 4820
rect 64230 4700 64236 4752
rect 64288 4740 64294 4752
rect 64325 4743 64383 4749
rect 64325 4740 64337 4743
rect 64288 4712 64337 4740
rect 64288 4700 64294 4712
rect 64325 4709 64337 4712
rect 64371 4709 64383 4743
rect 65610 4740 65616 4752
rect 65550 4712 65616 4740
rect 64325 4703 64383 4709
rect 65610 4700 65616 4712
rect 65668 4700 65674 4752
rect 64046 4632 64052 4684
rect 64104 4632 64110 4684
rect 63572 4378 66424 4400
rect 63572 4326 64338 4378
rect 64390 4326 64402 4378
rect 64454 4326 64466 4378
rect 64518 4326 64530 4378
rect 64582 4326 64594 4378
rect 64646 4326 66424 4378
rect 63572 4304 66424 4326
rect 63402 4224 63408 4276
rect 63460 4264 63466 4276
rect 64230 4264 64236 4276
rect 63460 4236 64236 4264
rect 63460 4224 63466 4236
rect 64230 4224 64236 4236
rect 64288 4224 64294 4276
rect 63865 4063 63923 4069
rect 63865 4029 63877 4063
rect 63911 4029 63923 4063
rect 63865 4023 63923 4029
rect 63880 3992 63908 4023
rect 64046 3992 64052 4004
rect 63880 3964 64052 3992
rect 64046 3952 64052 3964
rect 64104 3952 64110 4004
rect 64138 3952 64144 4004
rect 64196 3952 64202 4004
rect 65150 3952 65156 4004
rect 65208 3952 65214 4004
rect 65613 3927 65671 3933
rect 65613 3893 65625 3927
rect 65659 3924 65671 3927
rect 65978 3924 65984 3936
rect 65659 3896 65984 3924
rect 65659 3893 65671 3896
rect 65613 3887 65671 3893
rect 65978 3884 65984 3896
rect 66036 3884 66042 3936
rect 63572 3834 66424 3856
rect 63572 3782 65258 3834
rect 65310 3782 65322 3834
rect 65374 3782 65386 3834
rect 65438 3782 65450 3834
rect 65502 3782 65514 3834
rect 65566 3782 66424 3834
rect 63572 3760 66424 3782
rect 64138 3680 64144 3732
rect 64196 3720 64202 3732
rect 64693 3723 64751 3729
rect 64693 3720 64705 3723
rect 64196 3692 64705 3720
rect 64196 3680 64202 3692
rect 64693 3689 64705 3692
rect 64739 3689 64751 3723
rect 64693 3683 64751 3689
rect 64230 3612 64236 3664
rect 64288 3612 64294 3664
rect 65061 3655 65119 3661
rect 65061 3621 65073 3655
rect 65107 3652 65119 3655
rect 65150 3652 65156 3664
rect 65107 3624 65156 3652
rect 65107 3621 65119 3624
rect 65061 3615 65119 3621
rect 65150 3612 65156 3624
rect 65208 3612 65214 3664
rect 63954 3476 63960 3528
rect 64012 3476 64018 3528
rect 64141 3519 64199 3525
rect 64141 3485 64153 3519
rect 64187 3516 64199 3519
rect 64187 3488 64920 3516
rect 64187 3485 64199 3488
rect 64141 3479 64199 3485
rect 64601 3451 64659 3457
rect 64601 3417 64613 3451
rect 64647 3448 64659 3451
rect 64690 3448 64696 3460
rect 64647 3420 64696 3448
rect 64647 3417 64659 3420
rect 64601 3411 64659 3417
rect 64690 3408 64696 3420
rect 64748 3408 64754 3460
rect 64892 3448 64920 3488
rect 64966 3476 64972 3528
rect 65024 3516 65030 3528
rect 65153 3519 65211 3525
rect 65153 3516 65165 3519
rect 65024 3488 65165 3516
rect 65024 3476 65030 3488
rect 65153 3485 65165 3488
rect 65199 3485 65211 3519
rect 65153 3479 65211 3485
rect 65337 3519 65395 3525
rect 65337 3485 65349 3519
rect 65383 3516 65395 3519
rect 66438 3516 66444 3528
rect 65383 3488 66444 3516
rect 65383 3485 65395 3488
rect 65337 3479 65395 3485
rect 66438 3476 66444 3488
rect 66496 3476 66502 3528
rect 65978 3448 65984 3460
rect 64892 3420 65984 3448
rect 65978 3408 65984 3420
rect 66036 3408 66042 3460
rect 63770 3340 63776 3392
rect 63828 3380 63834 3392
rect 64782 3380 64788 3392
rect 63828 3352 64788 3380
rect 63828 3340 63834 3352
rect 64782 3340 64788 3352
rect 64840 3340 64846 3392
rect 63572 3290 66424 3312
rect 63572 3238 64338 3290
rect 64390 3238 64402 3290
rect 64454 3238 64466 3290
rect 64518 3238 64530 3290
rect 64582 3238 64594 3290
rect 64646 3238 66424 3290
rect 63572 3216 66424 3238
rect 63957 3179 64015 3185
rect 63957 3145 63969 3179
rect 64003 3176 64015 3179
rect 64138 3176 64144 3188
rect 64003 3148 64144 3176
rect 64003 3145 64015 3148
rect 63957 3139 64015 3145
rect 64138 3136 64144 3148
rect 64196 3136 64202 3188
rect 64046 3000 64052 3052
rect 64104 3000 64110 3052
rect 65794 3000 65800 3052
rect 65852 3000 65858 3052
rect 64322 2864 64328 2916
rect 64380 2864 64386 2916
rect 65610 2904 65616 2916
rect 65550 2876 65616 2904
rect 65610 2864 65616 2876
rect 65668 2864 65674 2916
rect 63572 2746 66424 2768
rect 63572 2694 65258 2746
rect 65310 2694 65322 2746
rect 65374 2694 65386 2746
rect 65438 2694 65450 2746
rect 65502 2694 65514 2746
rect 65566 2694 66424 2746
rect 63572 2672 66424 2694
rect 64322 2592 64328 2644
rect 64380 2632 64386 2644
rect 64601 2635 64659 2641
rect 64601 2632 64613 2635
rect 64380 2604 64613 2632
rect 64380 2592 64386 2604
rect 64601 2601 64613 2604
rect 64647 2601 64659 2635
rect 64601 2595 64659 2601
rect 65153 2635 65211 2641
rect 65153 2601 65165 2635
rect 65199 2632 65211 2635
rect 65702 2632 65708 2644
rect 65199 2604 65708 2632
rect 65199 2601 65211 2604
rect 65153 2595 65211 2601
rect 65702 2592 65708 2604
rect 65760 2592 65766 2644
rect 65061 2567 65119 2573
rect 65061 2533 65073 2567
rect 65107 2564 65119 2567
rect 66346 2564 66352 2576
rect 65107 2536 66352 2564
rect 65107 2533 65119 2536
rect 65061 2527 65119 2533
rect 66346 2524 66352 2536
rect 66404 2524 66410 2576
rect 64233 2499 64291 2505
rect 64233 2465 64245 2499
rect 64279 2496 64291 2499
rect 64966 2496 64972 2508
rect 64279 2468 64972 2496
rect 64279 2465 64291 2468
rect 64233 2459 64291 2465
rect 64966 2456 64972 2468
rect 65024 2456 65030 2508
rect 64049 2431 64107 2437
rect 64049 2397 64061 2431
rect 64095 2397 64107 2431
rect 64049 2391 64107 2397
rect 64141 2431 64199 2437
rect 64141 2397 64153 2431
rect 64187 2428 64199 2431
rect 64187 2400 64736 2428
rect 64187 2397 64199 2400
rect 64141 2391 64199 2397
rect 64064 2292 64092 2391
rect 64708 2369 64736 2400
rect 64782 2388 64788 2440
rect 64840 2428 64846 2440
rect 65242 2428 65248 2440
rect 64840 2400 65248 2428
rect 64840 2388 64846 2400
rect 65242 2388 65248 2400
rect 65300 2388 65306 2440
rect 64693 2363 64751 2369
rect 64693 2329 64705 2363
rect 64739 2329 64751 2363
rect 64693 2323 64751 2329
rect 64874 2292 64880 2304
rect 64064 2264 64880 2292
rect 64874 2252 64880 2264
rect 64932 2252 64938 2304
rect 63572 2202 66424 2224
rect 63572 2150 64338 2202
rect 64390 2150 64402 2202
rect 64454 2150 64466 2202
rect 64518 2150 64530 2202
rect 64582 2150 64594 2202
rect 64646 2150 66424 2202
rect 63572 2128 66424 2150
rect 65058 2048 65064 2100
rect 65116 2088 65122 2100
rect 65429 2091 65487 2097
rect 65429 2088 65441 2091
rect 65116 2060 65441 2088
rect 65116 2048 65122 2060
rect 65429 2057 65441 2060
rect 65475 2057 65487 2091
rect 65429 2051 65487 2057
rect 49234 1980 49240 2032
rect 49292 2020 49298 2032
rect 62758 2020 62764 2032
rect 49292 1992 62764 2020
rect 49292 1980 49298 1992
rect 62758 1980 62764 1992
rect 62816 1980 62822 2032
rect 64601 2023 64659 2029
rect 64601 1989 64613 2023
rect 64647 2020 64659 2023
rect 66162 2020 66168 2032
rect 64647 1992 66168 2020
rect 64647 1989 64659 1992
rect 64601 1983 64659 1989
rect 66162 1980 66168 1992
rect 66220 1980 66226 2032
rect 48958 1912 48964 1964
rect 49016 1952 49022 1964
rect 62666 1952 62672 1964
rect 49016 1924 62672 1952
rect 49016 1912 49022 1924
rect 62666 1912 62672 1924
rect 62724 1912 62730 1964
rect 65242 1912 65248 1964
rect 65300 1912 65306 1964
rect 65702 1912 65708 1964
rect 65760 1952 65766 1964
rect 65981 1955 66039 1961
rect 65981 1952 65993 1955
rect 65760 1924 65993 1952
rect 65760 1912 65766 1924
rect 65981 1921 65993 1924
rect 66027 1921 66039 1955
rect 65981 1915 66039 1921
rect 49694 1844 49700 1896
rect 49752 1884 49758 1896
rect 63034 1884 63040 1896
rect 49752 1856 63040 1884
rect 49752 1844 49758 1856
rect 63034 1844 63040 1856
rect 63092 1844 63098 1896
rect 64690 1844 64696 1896
rect 64748 1884 64754 1896
rect 64969 1887 65027 1893
rect 64969 1884 64981 1887
rect 64748 1856 64981 1884
rect 64748 1844 64754 1856
rect 64969 1853 64981 1856
rect 65015 1853 65027 1887
rect 64969 1847 65027 1853
rect 65061 1887 65119 1893
rect 65061 1853 65073 1887
rect 65107 1884 65119 1887
rect 65794 1884 65800 1896
rect 65107 1856 65800 1884
rect 65107 1853 65119 1856
rect 65061 1847 65119 1853
rect 65794 1844 65800 1856
rect 65852 1844 65858 1896
rect 63572 1658 66424 1680
rect 63572 1606 65258 1658
rect 65310 1606 65322 1658
rect 65374 1606 65386 1658
rect 65438 1606 65450 1658
rect 65502 1606 65514 1658
rect 65566 1606 66424 1658
rect 63572 1584 66424 1606
rect 65150 1504 65156 1556
rect 65208 1544 65214 1556
rect 65429 1547 65487 1553
rect 65429 1544 65441 1547
rect 65208 1516 65441 1544
rect 65208 1504 65214 1516
rect 65429 1513 65441 1516
rect 65475 1513 65487 1547
rect 65429 1507 65487 1513
rect 64690 1300 64696 1352
rect 64748 1300 64754 1352
rect 65978 1300 65984 1352
rect 66036 1300 66042 1352
rect 63572 1114 66424 1136
rect 63572 1062 64338 1114
rect 64390 1062 64402 1114
rect 64454 1062 64466 1114
rect 64518 1062 64530 1114
rect 64582 1062 64594 1114
rect 64646 1062 66424 1114
rect 63572 1040 66424 1062
rect 64966 960 64972 1012
rect 65024 1000 65030 1012
rect 65429 1003 65487 1009
rect 65429 1000 65441 1003
rect 65024 972 65441 1000
rect 65024 960 65030 972
rect 65429 969 65441 972
rect 65475 969 65487 1003
rect 65429 963 65487 969
rect 65794 824 65800 876
rect 65852 864 65858 876
rect 65981 867 66039 873
rect 65981 864 65993 867
rect 65852 836 65993 864
rect 65852 824 65858 836
rect 65981 833 65993 836
rect 66027 833 66039 867
rect 65981 827 66039 833
rect 63572 570 66424 592
rect 63572 518 65258 570
rect 65310 518 65322 570
rect 65374 518 65386 570
rect 65438 518 65450 570
rect 65502 518 65514 570
rect 65566 518 66424 570
rect 63572 496 66424 518
<< via1 >>
rect 27712 44820 27764 44872
rect 28816 44820 28868 44872
rect 30932 44820 30984 44872
rect 16764 44752 16816 44804
rect 21732 44752 21784 44804
rect 24860 44752 24912 44804
rect 33508 44752 33560 44804
rect 17316 44684 17368 44736
rect 24032 44684 24084 44736
rect 29184 44684 29236 44736
rect 40408 44684 40460 44736
rect 1998 44582 2050 44634
rect 2062 44582 2114 44634
rect 2126 44582 2178 44634
rect 2190 44582 2242 44634
rect 2254 44582 2306 44634
rect 50998 44582 51050 44634
rect 51062 44582 51114 44634
rect 51126 44582 51178 44634
rect 51190 44582 51242 44634
rect 51254 44582 51306 44634
rect 6184 44523 6236 44532
rect 6184 44489 6193 44523
rect 6193 44489 6227 44523
rect 6227 44489 6236 44523
rect 6184 44480 6236 44489
rect 6736 44523 6788 44532
rect 6736 44489 6745 44523
rect 6745 44489 6779 44523
rect 6779 44489 6788 44523
rect 6736 44480 6788 44489
rect 7288 44523 7340 44532
rect 7288 44489 7297 44523
rect 7297 44489 7331 44523
rect 7331 44489 7340 44523
rect 7288 44480 7340 44489
rect 7840 44523 7892 44532
rect 7840 44489 7849 44523
rect 7849 44489 7883 44523
rect 7883 44489 7892 44523
rect 7840 44480 7892 44489
rect 8392 44523 8444 44532
rect 8392 44489 8401 44523
rect 8401 44489 8435 44523
rect 8435 44489 8444 44523
rect 8392 44480 8444 44489
rect 8944 44523 8996 44532
rect 8944 44489 8953 44523
rect 8953 44489 8987 44523
rect 8987 44489 8996 44523
rect 8944 44480 8996 44489
rect 9496 44523 9548 44532
rect 9496 44489 9505 44523
rect 9505 44489 9539 44523
rect 9539 44489 9548 44523
rect 9496 44480 9548 44489
rect 10048 44523 10100 44532
rect 10048 44489 10057 44523
rect 10057 44489 10091 44523
rect 10091 44489 10100 44523
rect 10048 44480 10100 44489
rect 10600 44523 10652 44532
rect 10600 44489 10609 44523
rect 10609 44489 10643 44523
rect 10643 44489 10652 44523
rect 10600 44480 10652 44489
rect 12256 44523 12308 44532
rect 12256 44489 12265 44523
rect 12265 44489 12299 44523
rect 12299 44489 12308 44523
rect 12256 44480 12308 44489
rect 12532 44523 12584 44532
rect 12532 44489 12541 44523
rect 12541 44489 12575 44523
rect 12575 44489 12584 44523
rect 12532 44480 12584 44489
rect 12808 44523 12860 44532
rect 12808 44489 12817 44523
rect 12817 44489 12851 44523
rect 12851 44489 12860 44523
rect 12808 44480 12860 44489
rect 13544 44523 13596 44532
rect 13544 44489 13553 44523
rect 13553 44489 13587 44523
rect 13587 44489 13596 44523
rect 13544 44480 13596 44489
rect 13820 44523 13872 44532
rect 13820 44489 13829 44523
rect 13829 44489 13863 44523
rect 13863 44489 13872 44523
rect 13820 44480 13872 44489
rect 15476 44523 15528 44532
rect 15476 44489 15485 44523
rect 15485 44489 15519 44523
rect 15519 44489 15528 44523
rect 15476 44480 15528 44489
rect 15936 44523 15988 44532
rect 15936 44489 15945 44523
rect 15945 44489 15979 44523
rect 15979 44489 15988 44523
rect 15936 44480 15988 44489
rect 16212 44523 16264 44532
rect 16212 44489 16221 44523
rect 16221 44489 16255 44523
rect 16255 44489 16264 44523
rect 16212 44480 16264 44489
rect 16672 44523 16724 44532
rect 16672 44489 16681 44523
rect 16681 44489 16715 44523
rect 16715 44489 16724 44523
rect 16672 44480 16724 44489
rect 16948 44523 17000 44532
rect 16948 44489 16957 44523
rect 16957 44489 16991 44523
rect 16991 44489 17000 44523
rect 16948 44480 17000 44489
rect 17224 44523 17276 44532
rect 17224 44489 17233 44523
rect 17233 44489 17267 44523
rect 17267 44489 17276 44523
rect 17224 44480 17276 44489
rect 20076 44480 20128 44532
rect 21732 44480 21784 44532
rect 12256 44276 12308 44328
rect 14372 44276 14424 44328
rect 26424 44412 26476 44464
rect 17868 44344 17920 44396
rect 18512 44319 18564 44328
rect 18512 44285 18521 44319
rect 18521 44285 18555 44319
rect 18555 44285 18564 44319
rect 18512 44276 18564 44285
rect 19156 44276 19208 44328
rect 10600 44208 10652 44260
rect 11612 44183 11664 44192
rect 11612 44149 11621 44183
rect 11621 44149 11655 44183
rect 11655 44149 11664 44183
rect 11612 44140 11664 44149
rect 14188 44208 14240 44260
rect 18880 44208 18932 44260
rect 22284 44344 22336 44396
rect 20720 44208 20772 44260
rect 20996 44208 21048 44260
rect 21456 44208 21508 44260
rect 23940 44344 23992 44396
rect 22560 44276 22612 44328
rect 24032 44319 24084 44328
rect 24032 44285 24041 44319
rect 24041 44285 24075 44319
rect 24075 44285 24084 44319
rect 24032 44276 24084 44285
rect 26240 44276 26292 44328
rect 26608 44319 26660 44328
rect 26608 44285 26617 44319
rect 26617 44285 26651 44319
rect 26651 44285 26660 44319
rect 26608 44276 26660 44285
rect 26792 44387 26844 44396
rect 26792 44353 26801 44387
rect 26801 44353 26835 44387
rect 26835 44353 26844 44387
rect 26792 44344 26844 44353
rect 27528 44387 27580 44396
rect 27528 44353 27537 44387
rect 27537 44353 27571 44387
rect 27571 44353 27580 44387
rect 27528 44344 27580 44353
rect 27436 44276 27488 44328
rect 28632 44276 28684 44328
rect 30472 44276 30524 44328
rect 30932 44480 30984 44532
rect 36544 44480 36596 44532
rect 33048 44344 33100 44396
rect 35716 44344 35768 44396
rect 31852 44276 31904 44328
rect 34244 44276 34296 44328
rect 35440 44276 35492 44328
rect 38108 44412 38160 44464
rect 37924 44344 37976 44396
rect 38016 44387 38068 44396
rect 38016 44353 38025 44387
rect 38025 44353 38059 44387
rect 38059 44353 38068 44387
rect 38016 44344 38068 44353
rect 41604 44480 41656 44532
rect 42524 44480 42576 44532
rect 38292 44412 38344 44464
rect 39396 44412 39448 44464
rect 38292 44319 38344 44328
rect 38292 44285 38301 44319
rect 38301 44285 38335 44319
rect 38335 44285 38344 44319
rect 38292 44276 38344 44285
rect 39856 44276 39908 44328
rect 40408 44319 40460 44328
rect 40408 44285 40417 44319
rect 40417 44285 40451 44319
rect 40451 44285 40460 44319
rect 40408 44276 40460 44285
rect 42524 44387 42576 44396
rect 42524 44353 42533 44387
rect 42533 44353 42567 44387
rect 42567 44353 42576 44387
rect 42524 44344 42576 44353
rect 43076 44344 43128 44396
rect 43996 44344 44048 44396
rect 23388 44208 23440 44260
rect 26056 44251 26108 44260
rect 26056 44217 26065 44251
rect 26065 44217 26099 44251
rect 26099 44217 26108 44251
rect 26056 44208 26108 44217
rect 12532 44140 12584 44192
rect 12900 44140 12952 44192
rect 14740 44140 14792 44192
rect 14832 44140 14884 44192
rect 17500 44140 17552 44192
rect 17592 44140 17644 44192
rect 18972 44140 19024 44192
rect 20260 44140 20312 44192
rect 21548 44140 21600 44192
rect 22100 44140 22152 44192
rect 22468 44140 22520 44192
rect 25044 44183 25096 44192
rect 25044 44149 25053 44183
rect 25053 44149 25087 44183
rect 25087 44149 25096 44183
rect 25044 44140 25096 44149
rect 25320 44140 25372 44192
rect 25504 44183 25556 44192
rect 25504 44149 25513 44183
rect 25513 44149 25547 44183
rect 25547 44149 25556 44183
rect 25504 44140 25556 44149
rect 25596 44140 25648 44192
rect 27344 44183 27396 44192
rect 27344 44149 27353 44183
rect 27353 44149 27387 44183
rect 27387 44149 27396 44183
rect 27344 44140 27396 44149
rect 28724 44140 28776 44192
rect 29184 44251 29236 44260
rect 29184 44217 29193 44251
rect 29193 44217 29227 44251
rect 29227 44217 29236 44251
rect 29184 44208 29236 44217
rect 30840 44208 30892 44260
rect 29368 44183 29420 44192
rect 29368 44149 29377 44183
rect 29377 44149 29411 44183
rect 29411 44149 29420 44183
rect 29368 44140 29420 44149
rect 30748 44140 30800 44192
rect 32404 44140 32456 44192
rect 33324 44183 33376 44192
rect 33324 44149 33333 44183
rect 33333 44149 33367 44183
rect 33367 44149 33376 44183
rect 33324 44140 33376 44149
rect 33416 44183 33468 44192
rect 33416 44149 33425 44183
rect 33425 44149 33459 44183
rect 33459 44149 33468 44183
rect 33416 44140 33468 44149
rect 33968 44140 34020 44192
rect 35532 44140 35584 44192
rect 36636 44140 36688 44192
rect 37464 44183 37516 44192
rect 37464 44149 37473 44183
rect 37473 44149 37507 44183
rect 37507 44149 37516 44183
rect 37464 44140 37516 44149
rect 37740 44208 37792 44260
rect 38108 44208 38160 44260
rect 38752 44208 38804 44260
rect 38844 44140 38896 44192
rect 39028 44140 39080 44192
rect 39580 44140 39632 44192
rect 40500 44208 40552 44260
rect 40868 44208 40920 44260
rect 43812 44276 43864 44328
rect 48228 44344 48280 44396
rect 47400 44276 47452 44328
rect 50344 44208 50396 44260
rect 41512 44140 41564 44192
rect 42248 44183 42300 44192
rect 42248 44149 42257 44183
rect 42257 44149 42291 44183
rect 42291 44149 42300 44183
rect 42248 44140 42300 44149
rect 42340 44183 42392 44192
rect 42340 44149 42349 44183
rect 42349 44149 42383 44183
rect 42383 44149 42392 44183
rect 42340 44140 42392 44149
rect 42432 44140 42484 44192
rect 44456 44140 44508 44192
rect 45376 44140 45428 44192
rect 46940 44140 46992 44192
rect 2918 44038 2970 44090
rect 2982 44038 3034 44090
rect 3046 44038 3098 44090
rect 3110 44038 3162 44090
rect 3174 44038 3226 44090
rect 51918 44038 51970 44090
rect 51982 44038 52034 44090
rect 52046 44038 52098 44090
rect 52110 44038 52162 44090
rect 52174 44038 52226 44090
rect 11612 43936 11664 43988
rect 14372 43979 14424 43988
rect 14372 43945 14381 43979
rect 14381 43945 14415 43979
rect 14415 43945 14424 43979
rect 14372 43936 14424 43945
rect 14832 43979 14884 43988
rect 14832 43945 14841 43979
rect 14841 43945 14875 43979
rect 14875 43945 14884 43979
rect 14832 43936 14884 43945
rect 16120 43936 16172 43988
rect 12992 43868 13044 43920
rect 16856 43868 16908 43920
rect 17316 43911 17368 43920
rect 17316 43877 17325 43911
rect 17325 43877 17359 43911
rect 17359 43877 17368 43911
rect 17316 43868 17368 43877
rect 17500 43868 17552 43920
rect 18972 43868 19024 43920
rect 24124 43936 24176 43988
rect 11152 43843 11204 43852
rect 11152 43809 11161 43843
rect 11161 43809 11195 43843
rect 11195 43809 11204 43843
rect 11152 43800 11204 43809
rect 12532 43800 12584 43852
rect 14740 43800 14792 43852
rect 12440 43732 12492 43784
rect 15292 43843 15344 43852
rect 15292 43809 15301 43843
rect 15301 43809 15335 43843
rect 15335 43809 15344 43843
rect 15292 43800 15344 43809
rect 15660 43843 15712 43852
rect 15660 43809 15669 43843
rect 15669 43809 15703 43843
rect 15703 43809 15712 43843
rect 15660 43800 15712 43809
rect 20720 43868 20772 43920
rect 21548 43911 21600 43920
rect 21548 43877 21557 43911
rect 21557 43877 21591 43911
rect 21591 43877 21600 43911
rect 21548 43868 21600 43877
rect 22192 43868 22244 43920
rect 24952 43868 25004 43920
rect 26240 43936 26292 43988
rect 26884 43936 26936 43988
rect 16396 43732 16448 43784
rect 19524 43800 19576 43852
rect 19800 43732 19852 43784
rect 19892 43775 19944 43784
rect 19892 43741 19901 43775
rect 19901 43741 19935 43775
rect 19935 43741 19944 43775
rect 19892 43732 19944 43741
rect 20628 43732 20680 43784
rect 20812 43843 20864 43852
rect 20812 43809 20821 43843
rect 20821 43809 20855 43843
rect 20855 43809 20864 43843
rect 20812 43800 20864 43809
rect 22836 43800 22888 43852
rect 23388 43800 23440 43852
rect 26240 43843 26292 43852
rect 26240 43809 26249 43843
rect 26249 43809 26283 43843
rect 26283 43809 26292 43843
rect 26240 43800 26292 43809
rect 27344 43911 27396 43920
rect 27344 43877 27353 43911
rect 27353 43877 27387 43911
rect 27387 43877 27396 43911
rect 27344 43868 27396 43877
rect 27712 43868 27764 43920
rect 28908 43800 28960 43852
rect 29644 43911 29696 43920
rect 29644 43877 29653 43911
rect 29653 43877 29687 43911
rect 29687 43877 29696 43911
rect 29644 43868 29696 43877
rect 30656 43800 30708 43852
rect 22284 43732 22336 43784
rect 22744 43732 22796 43784
rect 25320 43732 25372 43784
rect 25964 43775 26016 43784
rect 25964 43741 25973 43775
rect 25973 43741 26007 43775
rect 26007 43741 26016 43775
rect 25964 43732 26016 43741
rect 26332 43732 26384 43784
rect 27068 43732 27120 43784
rect 29000 43732 29052 43784
rect 30380 43732 30432 43784
rect 31392 43775 31444 43784
rect 31392 43741 31401 43775
rect 31401 43741 31435 43775
rect 31435 43741 31444 43775
rect 31392 43732 31444 43741
rect 11060 43596 11112 43648
rect 12716 43596 12768 43648
rect 14740 43596 14792 43648
rect 17960 43664 18012 43716
rect 24584 43664 24636 43716
rect 36636 43936 36688 43988
rect 37280 43936 37332 43988
rect 38292 43936 38344 43988
rect 38844 43936 38896 43988
rect 41052 43936 41104 43988
rect 42248 43936 42300 43988
rect 47400 43979 47452 43988
rect 47400 43945 47409 43979
rect 47409 43945 47443 43979
rect 47443 43945 47452 43979
rect 47400 43936 47452 43945
rect 33968 43911 34020 43920
rect 33968 43877 33977 43911
rect 33977 43877 34011 43911
rect 34011 43877 34020 43911
rect 33968 43868 34020 43877
rect 34060 43868 34112 43920
rect 38108 43868 38160 43920
rect 38660 43868 38712 43920
rect 31852 43843 31904 43852
rect 31852 43809 31861 43843
rect 31861 43809 31895 43843
rect 31895 43809 31904 43843
rect 31852 43800 31904 43809
rect 36636 43800 36688 43852
rect 38936 43843 38988 43852
rect 38936 43809 38945 43843
rect 38945 43809 38979 43843
rect 38979 43809 38988 43843
rect 38936 43800 38988 43809
rect 39396 43843 39448 43852
rect 39396 43809 39405 43843
rect 39405 43809 39439 43843
rect 39439 43809 39448 43843
rect 39396 43800 39448 43809
rect 32220 43775 32272 43784
rect 32220 43741 32229 43775
rect 32229 43741 32263 43775
rect 32263 43741 32272 43775
rect 32220 43732 32272 43741
rect 33048 43775 33100 43784
rect 33048 43741 33057 43775
rect 33057 43741 33091 43775
rect 33091 43741 33100 43775
rect 33048 43732 33100 43741
rect 33600 43732 33652 43784
rect 18052 43596 18104 43648
rect 19248 43596 19300 43648
rect 19432 43639 19484 43648
rect 19432 43605 19441 43639
rect 19441 43605 19475 43639
rect 19475 43605 19484 43639
rect 19432 43596 19484 43605
rect 20076 43596 20128 43648
rect 21916 43596 21968 43648
rect 22652 43596 22704 43648
rect 26240 43596 26292 43648
rect 26516 43596 26568 43648
rect 32128 43664 32180 43716
rect 35440 43775 35492 43784
rect 35440 43741 35449 43775
rect 35449 43741 35483 43775
rect 35483 43741 35492 43775
rect 35440 43732 35492 43741
rect 35532 43707 35584 43716
rect 35532 43673 35541 43707
rect 35541 43673 35575 43707
rect 35575 43673 35584 43707
rect 35532 43664 35584 43673
rect 31668 43639 31720 43648
rect 31668 43605 31677 43639
rect 31677 43605 31711 43639
rect 31711 43605 31720 43639
rect 31668 43596 31720 43605
rect 33232 43596 33284 43648
rect 33692 43596 33744 43648
rect 34336 43596 34388 43648
rect 37556 43732 37608 43784
rect 42432 43868 42484 43920
rect 42892 43868 42944 43920
rect 45376 43911 45428 43920
rect 45376 43877 45385 43911
rect 45385 43877 45419 43911
rect 45419 43877 45428 43911
rect 45376 43868 45428 43877
rect 46020 43868 46072 43920
rect 39948 43800 40000 43852
rect 36636 43596 36688 43648
rect 40224 43732 40276 43784
rect 40776 43732 40828 43784
rect 39580 43707 39632 43716
rect 39580 43673 39589 43707
rect 39589 43673 39623 43707
rect 39623 43673 39632 43707
rect 39580 43664 39632 43673
rect 41972 43732 42024 43784
rect 42708 43732 42760 43784
rect 48044 43800 48096 43852
rect 43812 43775 43864 43784
rect 43812 43741 43821 43775
rect 43821 43741 43855 43775
rect 43855 43741 43864 43775
rect 43812 43732 43864 43741
rect 45100 43775 45152 43784
rect 45100 43741 45109 43775
rect 45109 43741 45143 43775
rect 45143 43741 45152 43775
rect 45100 43732 45152 43741
rect 47216 43732 47268 43784
rect 47584 43775 47636 43784
rect 47584 43741 47593 43775
rect 47593 43741 47627 43775
rect 47627 43741 47636 43775
rect 47584 43732 47636 43741
rect 48688 43775 48740 43784
rect 48688 43741 48697 43775
rect 48697 43741 48731 43775
rect 48731 43741 48740 43775
rect 48688 43732 48740 43741
rect 39304 43639 39356 43648
rect 39304 43605 39313 43639
rect 39313 43605 39347 43639
rect 39347 43605 39356 43639
rect 39304 43596 39356 43605
rect 41420 43596 41472 43648
rect 47308 43596 47360 43648
rect 47768 43596 47820 43648
rect 49424 43596 49476 43648
rect 1998 43494 2050 43546
rect 2062 43494 2114 43546
rect 2126 43494 2178 43546
rect 2190 43494 2242 43546
rect 2254 43494 2306 43546
rect 50998 43494 51050 43546
rect 51062 43494 51114 43546
rect 51126 43494 51178 43546
rect 51190 43494 51242 43546
rect 51254 43494 51306 43546
rect 11060 43299 11112 43308
rect 11060 43265 11069 43299
rect 11069 43265 11103 43299
rect 11103 43265 11112 43299
rect 11060 43256 11112 43265
rect 12716 43392 12768 43444
rect 14004 43392 14056 43444
rect 16856 43392 16908 43444
rect 16948 43392 17000 43444
rect 17500 43392 17552 43444
rect 19616 43392 19668 43444
rect 19892 43392 19944 43444
rect 18788 43367 18840 43376
rect 18788 43333 18797 43367
rect 18797 43333 18831 43367
rect 18831 43333 18840 43367
rect 18788 43324 18840 43333
rect 21916 43435 21968 43444
rect 21916 43401 21925 43435
rect 21925 43401 21959 43435
rect 21959 43401 21968 43435
rect 21916 43392 21968 43401
rect 22100 43435 22152 43444
rect 22100 43401 22109 43435
rect 22109 43401 22143 43435
rect 22143 43401 22152 43435
rect 22100 43392 22152 43401
rect 23940 43435 23992 43444
rect 23940 43401 23949 43435
rect 23949 43401 23983 43435
rect 23983 43401 23992 43435
rect 23940 43392 23992 43401
rect 23572 43324 23624 43376
rect 25596 43392 25648 43444
rect 25964 43392 26016 43444
rect 28632 43435 28684 43444
rect 28632 43401 28641 43435
rect 28641 43401 28675 43435
rect 28675 43401 28684 43435
rect 28632 43392 28684 43401
rect 29000 43435 29052 43444
rect 29000 43401 29009 43435
rect 29009 43401 29043 43435
rect 29043 43401 29052 43435
rect 29000 43392 29052 43401
rect 29644 43392 29696 43444
rect 30104 43392 30156 43444
rect 31576 43392 31628 43444
rect 33140 43392 33192 43444
rect 33324 43392 33376 43444
rect 34244 43392 34296 43444
rect 36544 43392 36596 43444
rect 36636 43435 36688 43444
rect 36636 43401 36645 43435
rect 36645 43401 36679 43435
rect 36679 43401 36688 43435
rect 36636 43392 36688 43401
rect 37924 43392 37976 43444
rect 40132 43392 40184 43444
rect 16120 43256 16172 43308
rect 19064 43256 19116 43308
rect 19340 43256 19392 43308
rect 19616 43256 19668 43308
rect 20168 43256 20220 43308
rect 20720 43256 20772 43308
rect 16028 43231 16080 43240
rect 16028 43197 16037 43231
rect 16037 43197 16071 43231
rect 16071 43197 16080 43231
rect 16028 43188 16080 43197
rect 16212 43231 16264 43240
rect 16212 43197 16221 43231
rect 16221 43197 16255 43231
rect 16255 43197 16264 43231
rect 16212 43188 16264 43197
rect 10600 43120 10652 43172
rect 11704 43163 11756 43172
rect 11704 43129 11713 43163
rect 11713 43129 11747 43163
rect 11747 43129 11756 43163
rect 11704 43120 11756 43129
rect 12992 43120 13044 43172
rect 12348 43052 12400 43104
rect 13176 43095 13228 43104
rect 13176 43061 13185 43095
rect 13185 43061 13219 43095
rect 13219 43061 13228 43095
rect 13176 43052 13228 43061
rect 13820 43163 13872 43172
rect 13820 43129 13829 43163
rect 13829 43129 13863 43163
rect 13863 43129 13872 43163
rect 13820 43120 13872 43129
rect 14280 43120 14332 43172
rect 16580 43120 16632 43172
rect 16948 43120 17000 43172
rect 19248 43188 19300 43240
rect 21732 43231 21784 43240
rect 21732 43197 21741 43231
rect 21741 43197 21775 43231
rect 21775 43197 21784 43231
rect 21732 43188 21784 43197
rect 15568 43052 15620 43104
rect 18512 43052 18564 43104
rect 19156 43052 19208 43104
rect 20076 43120 20128 43172
rect 22468 43256 22520 43308
rect 22652 43299 22704 43308
rect 22652 43265 22661 43299
rect 22661 43265 22695 43299
rect 22695 43265 22704 43299
rect 22652 43256 22704 43265
rect 25504 43324 25556 43376
rect 26240 43324 26292 43376
rect 26332 43324 26384 43376
rect 24584 43256 24636 43308
rect 22100 43120 22152 43172
rect 22008 43052 22060 43104
rect 22192 43052 22244 43104
rect 22928 43095 22980 43104
rect 22928 43061 22937 43095
rect 22937 43061 22971 43095
rect 22971 43061 22980 43095
rect 22928 43052 22980 43061
rect 23664 43188 23716 43240
rect 24124 43231 24176 43240
rect 24124 43197 24133 43231
rect 24133 43197 24167 43231
rect 24167 43197 24176 43231
rect 24124 43188 24176 43197
rect 23848 43120 23900 43172
rect 24584 43120 24636 43172
rect 24952 43120 25004 43172
rect 27620 43299 27672 43308
rect 27620 43265 27629 43299
rect 27629 43265 27663 43299
rect 27663 43265 27672 43299
rect 27620 43256 27672 43265
rect 28264 43324 28316 43376
rect 28908 43324 28960 43376
rect 30748 43324 30800 43376
rect 28356 43256 28408 43308
rect 29644 43299 29696 43308
rect 29644 43265 29653 43299
rect 29653 43265 29687 43299
rect 29687 43265 29696 43299
rect 29644 43256 29696 43265
rect 30104 43256 30156 43308
rect 33692 43299 33744 43308
rect 33692 43265 33701 43299
rect 33701 43265 33735 43299
rect 33735 43265 33744 43299
rect 33692 43256 33744 43265
rect 37096 43256 37148 43308
rect 37464 43299 37516 43308
rect 37464 43265 37473 43299
rect 37473 43265 37507 43299
rect 37507 43265 37516 43299
rect 37464 43256 37516 43265
rect 38936 43299 38988 43308
rect 38936 43265 38945 43299
rect 38945 43265 38979 43299
rect 38979 43265 38988 43299
rect 38936 43256 38988 43265
rect 40776 43256 40828 43308
rect 41328 43256 41380 43308
rect 42340 43392 42392 43444
rect 43076 43392 43128 43444
rect 42708 43367 42760 43376
rect 42708 43333 42717 43367
rect 42717 43333 42751 43367
rect 42751 43333 42760 43367
rect 42708 43324 42760 43333
rect 42616 43256 42668 43308
rect 43812 43324 43864 43376
rect 25136 43052 25188 43104
rect 25320 43052 25372 43104
rect 27252 43120 27304 43172
rect 28448 43231 28500 43240
rect 28448 43197 28457 43231
rect 28457 43197 28491 43231
rect 28491 43197 28500 43231
rect 28448 43188 28500 43197
rect 28724 43188 28776 43240
rect 29368 43231 29420 43240
rect 29368 43197 29377 43231
rect 29377 43197 29411 43231
rect 29411 43197 29420 43231
rect 29368 43188 29420 43197
rect 30564 43188 30616 43240
rect 31208 43231 31260 43240
rect 31208 43197 31217 43231
rect 31217 43197 31251 43231
rect 31251 43197 31260 43231
rect 31208 43188 31260 43197
rect 31576 43231 31628 43240
rect 31576 43197 31585 43231
rect 31585 43197 31619 43231
rect 31619 43197 31628 43231
rect 31576 43188 31628 43197
rect 34612 43188 34664 43240
rect 39764 43188 39816 43240
rect 40868 43231 40920 43240
rect 40868 43197 40877 43231
rect 40877 43197 40911 43231
rect 40911 43197 40920 43231
rect 40868 43188 40920 43197
rect 42892 43188 42944 43240
rect 43904 43188 43956 43240
rect 47216 43256 47268 43308
rect 47308 43299 47360 43308
rect 47308 43265 47317 43299
rect 47317 43265 47351 43299
rect 47351 43265 47360 43299
rect 47308 43256 47360 43265
rect 48688 43256 48740 43308
rect 28632 43120 28684 43172
rect 30196 43163 30248 43172
rect 30196 43129 30205 43163
rect 30205 43129 30239 43163
rect 30239 43129 30248 43163
rect 30196 43120 30248 43129
rect 31392 43120 31444 43172
rect 33232 43120 33284 43172
rect 33692 43120 33744 43172
rect 34060 43120 34112 43172
rect 26148 43052 26200 43104
rect 26516 43095 26568 43104
rect 26516 43061 26525 43095
rect 26525 43061 26559 43095
rect 26559 43061 26568 43095
rect 26516 43052 26568 43061
rect 27344 43052 27396 43104
rect 27436 43052 27488 43104
rect 29092 43052 29144 43104
rect 29736 43052 29788 43104
rect 30288 43095 30340 43104
rect 30288 43061 30297 43095
rect 30297 43061 30331 43095
rect 30331 43061 30340 43095
rect 30288 43052 30340 43061
rect 30564 43052 30616 43104
rect 32220 43095 32272 43104
rect 32220 43061 32229 43095
rect 32229 43061 32263 43095
rect 32263 43061 32272 43095
rect 32220 43052 32272 43061
rect 34336 43052 34388 43104
rect 35164 43163 35216 43172
rect 35164 43129 35173 43163
rect 35173 43129 35207 43163
rect 35207 43129 35216 43163
rect 35164 43120 35216 43129
rect 38752 43120 38804 43172
rect 40408 43163 40460 43172
rect 40408 43129 40417 43163
rect 40417 43129 40451 43163
rect 40451 43129 40460 43163
rect 40408 43120 40460 43129
rect 41512 43120 41564 43172
rect 39948 43052 40000 43104
rect 41052 43052 41104 43104
rect 43076 43052 43128 43104
rect 46020 43120 46072 43172
rect 47400 43120 47452 43172
rect 49976 43188 50028 43240
rect 51724 43188 51776 43240
rect 48136 43120 48188 43172
rect 49148 43163 49200 43172
rect 49148 43129 49157 43163
rect 49157 43129 49191 43163
rect 49191 43129 49200 43163
rect 49148 43120 49200 43129
rect 52368 43163 52420 43172
rect 52368 43129 52377 43163
rect 52377 43129 52411 43163
rect 52411 43129 52420 43163
rect 52368 43120 52420 43129
rect 43444 43052 43496 43104
rect 44916 43095 44968 43104
rect 44916 43061 44925 43095
rect 44925 43061 44959 43095
rect 44959 43061 44968 43095
rect 44916 43052 44968 43061
rect 51540 43052 51592 43104
rect 51816 43052 51868 43104
rect 2918 42950 2970 43002
rect 2982 42950 3034 43002
rect 3046 42950 3098 43002
rect 3110 42950 3162 43002
rect 3174 42950 3226 43002
rect 51918 42950 51970 43002
rect 51982 42950 52034 43002
rect 52046 42950 52098 43002
rect 52110 42950 52162 43002
rect 52174 42950 52226 43002
rect 11704 42848 11756 42900
rect 12256 42848 12308 42900
rect 12532 42848 12584 42900
rect 14004 42848 14056 42900
rect 14372 42848 14424 42900
rect 14740 42848 14792 42900
rect 16212 42848 16264 42900
rect 14188 42780 14240 42832
rect 13176 42712 13228 42764
rect 14556 42712 14608 42764
rect 15016 42712 15068 42764
rect 16672 42780 16724 42832
rect 16948 42780 17000 42832
rect 16120 42755 16172 42764
rect 16120 42721 16129 42755
rect 16129 42721 16163 42755
rect 16163 42721 16172 42755
rect 16120 42712 16172 42721
rect 19524 42848 19576 42900
rect 19984 42848 20036 42900
rect 20260 42891 20312 42900
rect 20260 42857 20269 42891
rect 20269 42857 20303 42891
rect 20303 42857 20312 42891
rect 20260 42848 20312 42857
rect 20168 42780 20220 42832
rect 20812 42848 20864 42900
rect 22560 42848 22612 42900
rect 22744 42891 22796 42900
rect 22744 42857 22753 42891
rect 22753 42857 22787 42891
rect 22787 42857 22796 42891
rect 22744 42848 22796 42857
rect 24216 42848 24268 42900
rect 25412 42848 25464 42900
rect 26148 42848 26200 42900
rect 26516 42848 26568 42900
rect 27712 42848 27764 42900
rect 38568 42848 38620 42900
rect 38660 42891 38712 42900
rect 38660 42857 38669 42891
rect 38669 42857 38703 42891
rect 38703 42857 38712 42891
rect 38660 42848 38712 42857
rect 39028 42891 39080 42900
rect 39028 42857 39037 42891
rect 39037 42857 39071 42891
rect 39071 42857 39080 42891
rect 39028 42848 39080 42857
rect 39304 42848 39356 42900
rect 40408 42848 40460 42900
rect 40776 42848 40828 42900
rect 41052 42891 41104 42900
rect 41052 42857 41061 42891
rect 41061 42857 41095 42891
rect 41095 42857 41104 42891
rect 41052 42848 41104 42857
rect 41420 42891 41472 42900
rect 41420 42857 41429 42891
rect 41429 42857 41463 42891
rect 41463 42857 41472 42891
rect 41420 42848 41472 42857
rect 43812 42848 43864 42900
rect 44916 42848 44968 42900
rect 46020 42848 46072 42900
rect 46940 42848 46992 42900
rect 47216 42848 47268 42900
rect 48688 42848 48740 42900
rect 49148 42848 49200 42900
rect 49424 42891 49476 42900
rect 49424 42857 49433 42891
rect 49433 42857 49467 42891
rect 49467 42857 49476 42891
rect 49424 42848 49476 42857
rect 13084 42644 13136 42696
rect 13544 42687 13596 42696
rect 13544 42653 13553 42687
rect 13553 42653 13587 42687
rect 13587 42653 13596 42687
rect 13544 42644 13596 42653
rect 14004 42644 14056 42696
rect 14648 42644 14700 42696
rect 15384 42687 15436 42696
rect 15384 42653 15393 42687
rect 15393 42653 15427 42687
rect 15427 42653 15436 42687
rect 15384 42644 15436 42653
rect 16764 42644 16816 42696
rect 19432 42644 19484 42696
rect 22100 42780 22152 42832
rect 24952 42780 25004 42832
rect 27252 42823 27304 42832
rect 27252 42789 27261 42823
rect 27261 42789 27295 42823
rect 27295 42789 27304 42823
rect 27252 42780 27304 42789
rect 27344 42823 27396 42832
rect 27344 42789 27353 42823
rect 27353 42789 27387 42823
rect 27387 42789 27396 42823
rect 27344 42780 27396 42789
rect 29000 42780 29052 42832
rect 30196 42780 30248 42832
rect 30380 42780 30432 42832
rect 32404 42823 32456 42832
rect 32404 42789 32413 42823
rect 32413 42789 32447 42823
rect 32447 42789 32456 42823
rect 32404 42780 32456 42789
rect 33692 42780 33744 42832
rect 34152 42780 34204 42832
rect 34336 42823 34388 42832
rect 34336 42789 34345 42823
rect 34345 42789 34379 42823
rect 34379 42789 34388 42823
rect 34336 42780 34388 42789
rect 35532 42780 35584 42832
rect 39948 42780 40000 42832
rect 42892 42780 42944 42832
rect 51816 42780 51868 42832
rect 20904 42712 20956 42764
rect 22376 42712 22428 42764
rect 25872 42755 25924 42764
rect 25872 42721 25881 42755
rect 25881 42721 25915 42755
rect 25915 42721 25924 42755
rect 25872 42712 25924 42721
rect 26424 42755 26476 42764
rect 26424 42721 26433 42755
rect 26433 42721 26467 42755
rect 26467 42721 26476 42755
rect 26424 42712 26476 42721
rect 13820 42576 13872 42628
rect 15016 42619 15068 42628
rect 15016 42585 15025 42619
rect 15025 42585 15059 42619
rect 15059 42585 15068 42619
rect 15016 42576 15068 42585
rect 21456 42687 21508 42696
rect 21456 42653 21465 42687
rect 21465 42653 21499 42687
rect 21499 42653 21508 42687
rect 21456 42644 21508 42653
rect 22560 42644 22612 42696
rect 22836 42687 22888 42696
rect 22836 42653 22845 42687
rect 22845 42653 22879 42687
rect 22879 42653 22888 42687
rect 22836 42644 22888 42653
rect 14280 42508 14332 42560
rect 17132 42508 17184 42560
rect 17960 42508 18012 42560
rect 19248 42508 19300 42560
rect 20812 42508 20864 42560
rect 22376 42508 22428 42560
rect 23388 42687 23440 42696
rect 23388 42653 23397 42687
rect 23397 42653 23431 42687
rect 23431 42653 23440 42687
rect 23388 42644 23440 42653
rect 26056 42644 26108 42696
rect 28816 42755 28868 42764
rect 28816 42721 28825 42755
rect 28825 42721 28859 42755
rect 28859 42721 28868 42755
rect 28816 42712 28868 42721
rect 24676 42576 24728 42628
rect 26608 42619 26660 42628
rect 26608 42585 26617 42619
rect 26617 42585 26651 42619
rect 26651 42585 26660 42619
rect 26608 42576 26660 42585
rect 23480 42508 23532 42560
rect 26700 42508 26752 42560
rect 27620 42644 27672 42696
rect 28172 42687 28224 42696
rect 28172 42653 28181 42687
rect 28181 42653 28215 42687
rect 28215 42653 28224 42687
rect 28172 42644 28224 42653
rect 28356 42687 28408 42696
rect 28356 42653 28365 42687
rect 28365 42653 28399 42687
rect 28399 42653 28408 42687
rect 28356 42644 28408 42653
rect 28632 42644 28684 42696
rect 30472 42712 30524 42764
rect 35072 42712 35124 42764
rect 36636 42712 36688 42764
rect 36820 42755 36872 42764
rect 36820 42721 36829 42755
rect 36829 42721 36863 42755
rect 36863 42721 36872 42755
rect 36820 42712 36872 42721
rect 37280 42755 37332 42764
rect 37280 42721 37289 42755
rect 37289 42721 37323 42755
rect 37323 42721 37332 42755
rect 37280 42712 37332 42721
rect 39120 42712 39172 42764
rect 40500 42755 40552 42764
rect 40500 42721 40509 42755
rect 40509 42721 40543 42755
rect 40543 42721 40552 42755
rect 40500 42712 40552 42721
rect 41328 42712 41380 42764
rect 43720 42712 43772 42764
rect 46572 42712 46624 42764
rect 48136 42712 48188 42764
rect 48228 42712 48280 42764
rect 29092 42687 29144 42696
rect 29092 42653 29101 42687
rect 29101 42653 29135 42687
rect 29135 42653 29144 42687
rect 29092 42644 29144 42653
rect 32128 42687 32180 42696
rect 32128 42653 32137 42687
rect 32137 42653 32171 42687
rect 32171 42653 32180 42687
rect 32128 42644 32180 42653
rect 33692 42644 33744 42696
rect 34520 42687 34572 42696
rect 34520 42653 34529 42687
rect 34529 42653 34563 42687
rect 34563 42653 34572 42687
rect 34520 42644 34572 42653
rect 34980 42644 35032 42696
rect 27804 42576 27856 42628
rect 29184 42576 29236 42628
rect 29736 42619 29788 42628
rect 29736 42585 29745 42619
rect 29745 42585 29779 42619
rect 29779 42585 29788 42619
rect 29736 42576 29788 42585
rect 30288 42576 30340 42628
rect 33416 42576 33468 42628
rect 37556 42644 37608 42696
rect 38016 42644 38068 42696
rect 38384 42644 38436 42696
rect 37740 42619 37792 42628
rect 37740 42585 37749 42619
rect 37749 42585 37783 42619
rect 37783 42585 37792 42619
rect 37740 42576 37792 42585
rect 39304 42644 39356 42696
rect 42064 42644 42116 42696
rect 43444 42644 43496 42696
rect 44180 42687 44232 42696
rect 41604 42576 41656 42628
rect 30104 42508 30156 42560
rect 34612 42508 34664 42560
rect 35072 42508 35124 42560
rect 35716 42508 35768 42560
rect 35900 42551 35952 42560
rect 35900 42517 35909 42551
rect 35909 42517 35943 42551
rect 35943 42517 35952 42551
rect 35900 42508 35952 42517
rect 37832 42551 37884 42560
rect 37832 42517 37841 42551
rect 37841 42517 37875 42551
rect 37875 42517 37884 42551
rect 37832 42508 37884 42517
rect 40500 42508 40552 42560
rect 42524 42508 42576 42560
rect 42616 42508 42668 42560
rect 44180 42653 44189 42687
rect 44189 42653 44223 42687
rect 44223 42653 44232 42687
rect 44180 42644 44232 42653
rect 45652 42644 45704 42696
rect 46388 42644 46440 42696
rect 47492 42687 47544 42696
rect 47492 42653 47501 42687
rect 47501 42653 47535 42687
rect 47535 42653 47544 42687
rect 47492 42644 47544 42653
rect 47768 42644 47820 42696
rect 48688 42687 48740 42696
rect 48688 42653 48697 42687
rect 48697 42653 48731 42687
rect 48731 42653 48740 42687
rect 48688 42644 48740 42653
rect 47584 42576 47636 42628
rect 43904 42551 43956 42560
rect 43904 42517 43913 42551
rect 43913 42517 43947 42551
rect 43947 42517 43956 42551
rect 43904 42508 43956 42517
rect 44088 42508 44140 42560
rect 47676 42508 47728 42560
rect 48780 42508 48832 42560
rect 49516 42687 49568 42696
rect 49516 42653 49525 42687
rect 49525 42653 49559 42687
rect 49559 42653 49568 42687
rect 49516 42644 49568 42653
rect 49976 42755 50028 42764
rect 49976 42721 49985 42755
rect 49985 42721 50019 42755
rect 50019 42721 50028 42755
rect 49976 42712 50028 42721
rect 51632 42712 51684 42764
rect 60004 42712 60056 42764
rect 50252 42687 50304 42696
rect 50252 42653 50261 42687
rect 50261 42653 50295 42687
rect 50295 42653 50304 42687
rect 50252 42644 50304 42653
rect 50344 42644 50396 42696
rect 50804 42644 50856 42696
rect 54024 42644 54076 42696
rect 54116 42687 54168 42696
rect 54116 42653 54125 42687
rect 54125 42653 54159 42687
rect 54159 42653 54168 42687
rect 54116 42644 54168 42653
rect 52368 42619 52420 42628
rect 52368 42585 52377 42619
rect 52377 42585 52411 42619
rect 52411 42585 52420 42619
rect 52368 42576 52420 42585
rect 51724 42551 51776 42560
rect 51724 42517 51733 42551
rect 51733 42517 51767 42551
rect 51767 42517 51776 42551
rect 51724 42508 51776 42517
rect 53104 42508 53156 42560
rect 65800 42508 65852 42560
rect 1998 42406 2050 42458
rect 2062 42406 2114 42458
rect 2126 42406 2178 42458
rect 2190 42406 2242 42458
rect 2254 42406 2306 42458
rect 50998 42406 51050 42458
rect 51062 42406 51114 42458
rect 51126 42406 51178 42458
rect 51190 42406 51242 42458
rect 51254 42406 51306 42458
rect 10416 42304 10468 42356
rect 10600 42168 10652 42220
rect 10968 42168 11020 42220
rect 13544 42304 13596 42356
rect 15200 42304 15252 42356
rect 16028 42304 16080 42356
rect 16488 42347 16540 42356
rect 16488 42313 16497 42347
rect 16497 42313 16531 42347
rect 16531 42313 16540 42347
rect 16488 42304 16540 42313
rect 16764 42347 16816 42356
rect 16764 42313 16773 42347
rect 16773 42313 16807 42347
rect 16807 42313 16816 42347
rect 16764 42304 16816 42313
rect 20720 42304 20772 42356
rect 20812 42304 20864 42356
rect 22100 42304 22152 42356
rect 22652 42304 22704 42356
rect 14188 42168 14240 42220
rect 14740 42211 14792 42220
rect 14740 42177 14749 42211
rect 14749 42177 14783 42211
rect 14783 42177 14792 42211
rect 14740 42168 14792 42177
rect 16672 42168 16724 42220
rect 17868 42168 17920 42220
rect 18052 42211 18104 42220
rect 18052 42177 18061 42211
rect 18061 42177 18095 42211
rect 18095 42177 18104 42211
rect 18052 42168 18104 42177
rect 18420 42168 18472 42220
rect 7932 42100 7984 42152
rect 9772 42100 9824 42152
rect 17132 42143 17184 42152
rect 17132 42109 17141 42143
rect 17141 42109 17175 42143
rect 17175 42109 17184 42143
rect 17132 42100 17184 42109
rect 23112 42236 23164 42288
rect 23204 42236 23256 42288
rect 19156 42211 19208 42220
rect 19156 42177 19165 42211
rect 19165 42177 19199 42211
rect 19199 42177 19208 42211
rect 19156 42168 19208 42177
rect 19248 42211 19300 42220
rect 19248 42177 19257 42211
rect 19257 42177 19291 42211
rect 19291 42177 19300 42211
rect 19248 42168 19300 42177
rect 21824 42168 21876 42220
rect 22560 42168 22612 42220
rect 23020 42211 23072 42220
rect 23020 42177 23029 42211
rect 23029 42177 23063 42211
rect 23063 42177 23072 42211
rect 23020 42168 23072 42177
rect 24584 42304 24636 42356
rect 25136 42304 25188 42356
rect 24768 42236 24820 42288
rect 25044 42168 25096 42220
rect 25964 42168 26016 42220
rect 26240 42211 26292 42220
rect 26240 42177 26249 42211
rect 26249 42177 26283 42211
rect 26283 42177 26292 42211
rect 26240 42168 26292 42177
rect 15016 42075 15068 42084
rect 15016 42041 15025 42075
rect 15025 42041 15059 42075
rect 15059 42041 15068 42075
rect 15016 42032 15068 42041
rect 16304 42032 16356 42084
rect 16948 42032 17000 42084
rect 22928 42100 22980 42152
rect 24216 42143 24268 42152
rect 24216 42109 24225 42143
rect 24225 42109 24259 42143
rect 24259 42109 24268 42143
rect 24216 42100 24268 42109
rect 24584 42100 24636 42152
rect 26884 42211 26936 42220
rect 26884 42177 26893 42211
rect 26893 42177 26927 42211
rect 26927 42177 26936 42211
rect 26884 42168 26936 42177
rect 27620 42168 27672 42220
rect 28632 42347 28684 42356
rect 28632 42313 28641 42347
rect 28641 42313 28675 42347
rect 28675 42313 28684 42347
rect 28632 42304 28684 42313
rect 29000 42347 29052 42356
rect 29000 42313 29009 42347
rect 29009 42313 29043 42347
rect 29043 42313 29052 42347
rect 29000 42304 29052 42313
rect 33600 42304 33652 42356
rect 35072 42347 35124 42356
rect 35072 42313 35081 42347
rect 35081 42313 35115 42347
rect 35115 42313 35124 42347
rect 35072 42304 35124 42313
rect 35164 42304 35216 42356
rect 36820 42304 36872 42356
rect 28540 42236 28592 42288
rect 30840 42236 30892 42288
rect 32312 42168 32364 42220
rect 33140 42168 33192 42220
rect 33416 42211 33468 42220
rect 33416 42177 33425 42211
rect 33425 42177 33459 42211
rect 33459 42177 33468 42211
rect 33416 42168 33468 42177
rect 10692 42007 10744 42016
rect 10692 41973 10701 42007
rect 10701 41973 10735 42007
rect 10735 41973 10744 42007
rect 10692 41964 10744 41973
rect 17684 41964 17736 42016
rect 17960 42007 18012 42016
rect 17960 41973 17969 42007
rect 17969 41973 18003 42007
rect 18003 41973 18012 42007
rect 17960 41964 18012 41973
rect 20536 42032 20588 42084
rect 25780 42032 25832 42084
rect 28264 42100 28316 42152
rect 28632 42100 28684 42152
rect 30196 42100 30248 42152
rect 22376 42007 22428 42016
rect 22376 41973 22385 42007
rect 22385 41973 22419 42007
rect 22419 41973 22428 42007
rect 22376 41964 22428 41973
rect 23204 42007 23256 42016
rect 23204 41973 23213 42007
rect 23213 41973 23247 42007
rect 23247 41973 23256 42007
rect 23204 41964 23256 41973
rect 24124 41964 24176 42016
rect 24216 41964 24268 42016
rect 25412 41964 25464 42016
rect 25872 41964 25924 42016
rect 30656 42032 30708 42084
rect 30748 42075 30800 42084
rect 30748 42041 30757 42075
rect 30757 42041 30791 42075
rect 30791 42041 30800 42075
rect 30748 42032 30800 42041
rect 33692 42100 33744 42152
rect 34796 42236 34848 42288
rect 38936 42347 38988 42356
rect 38936 42313 38945 42347
rect 38945 42313 38979 42347
rect 38979 42313 38988 42347
rect 38936 42304 38988 42313
rect 39304 42304 39356 42356
rect 42064 42347 42116 42356
rect 42064 42313 42073 42347
rect 42073 42313 42107 42347
rect 42107 42313 42116 42347
rect 42064 42304 42116 42313
rect 34612 42211 34664 42220
rect 34612 42177 34621 42211
rect 34621 42177 34655 42211
rect 34655 42177 34664 42211
rect 34612 42168 34664 42177
rect 31852 42032 31904 42084
rect 30380 41964 30432 42016
rect 30472 41964 30524 42016
rect 32404 42032 32456 42084
rect 32220 41964 32272 42016
rect 33416 42032 33468 42084
rect 34244 42032 34296 42084
rect 34428 42100 34480 42152
rect 35716 42211 35768 42220
rect 35716 42177 35725 42211
rect 35725 42177 35759 42211
rect 35759 42177 35768 42211
rect 35716 42168 35768 42177
rect 35808 42211 35860 42220
rect 35808 42177 35817 42211
rect 35817 42177 35851 42211
rect 35851 42177 35860 42211
rect 35808 42168 35860 42177
rect 37832 42168 37884 42220
rect 35900 42100 35952 42152
rect 36268 42100 36320 42152
rect 40040 42100 40092 42152
rect 40868 42236 40920 42288
rect 41604 42168 41656 42220
rect 42432 42168 42484 42220
rect 42616 42211 42668 42220
rect 42616 42177 42625 42211
rect 42625 42177 42659 42211
rect 42659 42177 42668 42211
rect 42616 42168 42668 42177
rect 34980 42032 35032 42084
rect 38752 42032 38804 42084
rect 39396 42032 39448 42084
rect 41696 42143 41748 42152
rect 41696 42109 41705 42143
rect 41705 42109 41739 42143
rect 41739 42109 41748 42143
rect 41696 42100 41748 42109
rect 42708 42100 42760 42152
rect 43352 42236 43404 42288
rect 51632 42304 51684 42356
rect 51724 42304 51776 42356
rect 43904 42236 43956 42288
rect 43996 42211 44048 42220
rect 43996 42177 44005 42211
rect 44005 42177 44039 42211
rect 44039 42177 44048 42211
rect 43996 42168 44048 42177
rect 44088 42100 44140 42152
rect 44180 42100 44232 42152
rect 45468 42168 45520 42220
rect 46940 42168 46992 42220
rect 47400 42211 47452 42220
rect 47400 42177 47409 42211
rect 47409 42177 47443 42211
rect 47443 42177 47452 42211
rect 47400 42168 47452 42177
rect 47676 42211 47728 42220
rect 47676 42177 47685 42211
rect 47685 42177 47719 42211
rect 47719 42177 47728 42211
rect 47676 42168 47728 42177
rect 48688 42168 48740 42220
rect 49056 42168 49108 42220
rect 51356 42168 51408 42220
rect 53104 42143 53156 42152
rect 53104 42109 53113 42143
rect 53113 42109 53147 42143
rect 53147 42109 53156 42143
rect 53104 42100 53156 42109
rect 33232 42007 33284 42016
rect 33232 41973 33241 42007
rect 33241 41973 33275 42007
rect 33275 41973 33284 42007
rect 33232 41964 33284 41973
rect 33324 41964 33376 42016
rect 39304 42007 39356 42016
rect 39304 41973 39313 42007
rect 39313 41973 39347 42007
rect 39347 41973 39356 42007
rect 39304 41964 39356 41973
rect 39856 41964 39908 42016
rect 40316 41964 40368 42016
rect 41880 42075 41932 42084
rect 41880 42041 41889 42075
rect 41889 42041 41923 42075
rect 41923 42041 41932 42075
rect 41880 42032 41932 42041
rect 43444 42032 43496 42084
rect 43628 42032 43680 42084
rect 46020 42032 46072 42084
rect 47032 42075 47084 42084
rect 47032 42041 47041 42075
rect 47041 42041 47075 42075
rect 47075 42041 47084 42075
rect 47032 42032 47084 42041
rect 48136 42032 48188 42084
rect 50620 42075 50672 42084
rect 50620 42041 50629 42075
rect 50629 42041 50663 42075
rect 50663 42041 50672 42075
rect 50620 42032 50672 42041
rect 51816 42032 51868 42084
rect 54208 42211 54260 42220
rect 54208 42177 54217 42211
rect 54217 42177 54251 42211
rect 54251 42177 54260 42211
rect 54208 42168 54260 42177
rect 54024 42100 54076 42152
rect 63040 42100 63092 42152
rect 43076 41964 43128 42016
rect 44456 42007 44508 42016
rect 44456 41973 44465 42007
rect 44465 41973 44499 42007
rect 44499 41973 44508 42007
rect 44456 41964 44508 41973
rect 44824 42007 44876 42016
rect 44824 41973 44833 42007
rect 44833 41973 44867 42007
rect 44867 41973 44876 42007
rect 44824 41964 44876 41973
rect 45560 42007 45612 42016
rect 45560 41973 45569 42007
rect 45569 41973 45603 42007
rect 45603 41973 45612 42007
rect 45560 41964 45612 41973
rect 46848 41964 46900 42016
rect 46940 41964 46992 42016
rect 52276 41964 52328 42016
rect 52460 41964 52512 42016
rect 53196 42007 53248 42016
rect 53196 41973 53205 42007
rect 53205 41973 53239 42007
rect 53239 41973 53248 42007
rect 53196 41964 53248 41973
rect 54484 42032 54536 42084
rect 54024 42007 54076 42016
rect 54024 41973 54033 42007
rect 54033 41973 54067 42007
rect 54067 41973 54076 42007
rect 54024 41964 54076 41973
rect 54852 42007 54904 42016
rect 54852 41973 54861 42007
rect 54861 41973 54895 42007
rect 54895 41973 54904 42007
rect 54852 41964 54904 41973
rect 2918 41862 2970 41914
rect 2982 41862 3034 41914
rect 3046 41862 3098 41914
rect 3110 41862 3162 41914
rect 3174 41862 3226 41914
rect 51918 41862 51970 41914
rect 51982 41862 52034 41914
rect 52046 41862 52098 41914
rect 52110 41862 52162 41914
rect 52174 41862 52226 41914
rect 10416 41803 10468 41812
rect 10416 41769 10425 41803
rect 10425 41769 10459 41803
rect 10459 41769 10468 41803
rect 10416 41760 10468 41769
rect 15016 41760 15068 41812
rect 15568 41803 15620 41812
rect 15568 41769 15577 41803
rect 15577 41769 15611 41803
rect 15611 41769 15620 41803
rect 15568 41760 15620 41769
rect 16580 41760 16632 41812
rect 17592 41803 17644 41812
rect 17592 41769 17601 41803
rect 17601 41769 17635 41803
rect 17635 41769 17644 41803
rect 17592 41760 17644 41769
rect 17684 41803 17736 41812
rect 17684 41769 17693 41803
rect 17693 41769 17727 41803
rect 17727 41769 17736 41803
rect 17684 41760 17736 41769
rect 20720 41760 20772 41812
rect 9772 41692 9824 41744
rect 15384 41692 15436 41744
rect 17960 41692 18012 41744
rect 23480 41760 23532 41812
rect 23664 41760 23716 41812
rect 23848 41760 23900 41812
rect 11428 41624 11480 41676
rect 7932 41599 7984 41608
rect 7932 41565 7941 41599
rect 7941 41565 7975 41599
rect 7975 41565 7984 41599
rect 7932 41556 7984 41565
rect 8208 41599 8260 41608
rect 8208 41565 8217 41599
rect 8217 41565 8251 41599
rect 8251 41565 8260 41599
rect 8208 41556 8260 41565
rect 10416 41556 10468 41608
rect 11336 41556 11388 41608
rect 12624 41556 12676 41608
rect 12900 41599 12952 41608
rect 12900 41565 12909 41599
rect 12909 41565 12943 41599
rect 12943 41565 12952 41599
rect 12900 41556 12952 41565
rect 13820 41599 13872 41608
rect 13820 41565 13829 41599
rect 13829 41565 13863 41599
rect 13863 41565 13872 41599
rect 13820 41556 13872 41565
rect 10968 41488 11020 41540
rect 13176 41488 13228 41540
rect 16672 41624 16724 41676
rect 16764 41667 16816 41676
rect 16764 41633 16773 41667
rect 16773 41633 16807 41667
rect 16807 41633 16816 41667
rect 16764 41624 16816 41633
rect 22192 41692 22244 41744
rect 23388 41692 23440 41744
rect 16396 41556 16448 41608
rect 17868 41599 17920 41608
rect 17868 41565 17877 41599
rect 17877 41565 17911 41599
rect 17911 41565 17920 41599
rect 17868 41556 17920 41565
rect 18328 41556 18380 41608
rect 18880 41488 18932 41540
rect 20628 41556 20680 41608
rect 20996 41599 21048 41608
rect 20996 41565 21005 41599
rect 21005 41565 21039 41599
rect 21039 41565 21048 41599
rect 20996 41556 21048 41565
rect 21548 41599 21600 41608
rect 21548 41565 21557 41599
rect 21557 41565 21591 41599
rect 21591 41565 21600 41599
rect 21548 41556 21600 41565
rect 22836 41556 22888 41608
rect 24216 41692 24268 41744
rect 24860 41692 24912 41744
rect 25780 41760 25832 41812
rect 27068 41760 27120 41812
rect 27528 41760 27580 41812
rect 23848 41667 23900 41676
rect 23848 41633 23857 41667
rect 23857 41633 23891 41667
rect 23891 41633 23900 41667
rect 23848 41624 23900 41633
rect 26700 41735 26752 41744
rect 26700 41701 26709 41735
rect 26709 41701 26743 41735
rect 26743 41701 26752 41735
rect 26700 41692 26752 41701
rect 28172 41760 28224 41812
rect 30840 41692 30892 41744
rect 32220 41735 32272 41744
rect 32220 41701 32229 41735
rect 32229 41701 32263 41735
rect 32263 41701 32272 41735
rect 32220 41692 32272 41701
rect 33692 41803 33744 41812
rect 33692 41769 33701 41803
rect 33701 41769 33735 41803
rect 33735 41769 33744 41803
rect 33692 41760 33744 41769
rect 39304 41760 39356 41812
rect 40224 41760 40276 41812
rect 41696 41760 41748 41812
rect 42524 41760 42576 41812
rect 37004 41692 37056 41744
rect 37096 41692 37148 41744
rect 38568 41692 38620 41744
rect 26240 41624 26292 41676
rect 23756 41599 23808 41608
rect 23756 41565 23765 41599
rect 23765 41565 23799 41599
rect 23799 41565 23808 41599
rect 23756 41556 23808 41565
rect 24124 41599 24176 41608
rect 24124 41565 24133 41599
rect 24133 41565 24167 41599
rect 24167 41565 24176 41599
rect 24124 41556 24176 41565
rect 25136 41556 25188 41608
rect 28540 41624 28592 41676
rect 30104 41624 30156 41676
rect 33324 41624 33376 41676
rect 34060 41624 34112 41676
rect 34980 41624 35032 41676
rect 9680 41463 9732 41472
rect 9680 41429 9689 41463
rect 9689 41429 9723 41463
rect 9723 41429 9732 41463
rect 9680 41420 9732 41429
rect 10048 41463 10100 41472
rect 10048 41429 10057 41463
rect 10057 41429 10091 41463
rect 10091 41429 10100 41463
rect 10048 41420 10100 41429
rect 10784 41420 10836 41472
rect 11888 41420 11940 41472
rect 14648 41420 14700 41472
rect 15384 41420 15436 41472
rect 16396 41420 16448 41472
rect 18052 41463 18104 41472
rect 18052 41429 18061 41463
rect 18061 41429 18095 41463
rect 18095 41429 18104 41463
rect 18052 41420 18104 41429
rect 19616 41463 19668 41472
rect 19616 41429 19625 41463
rect 19625 41429 19659 41463
rect 19659 41429 19668 41463
rect 19616 41420 19668 41429
rect 20260 41420 20312 41472
rect 21272 41488 21324 41540
rect 25872 41488 25924 41540
rect 28448 41556 28500 41608
rect 29184 41599 29236 41608
rect 29184 41565 29193 41599
rect 29193 41565 29227 41599
rect 29227 41565 29236 41599
rect 29184 41556 29236 41565
rect 27712 41488 27764 41540
rect 30380 41531 30432 41540
rect 30380 41497 30389 41531
rect 30389 41497 30423 41531
rect 30423 41497 30432 41531
rect 30380 41488 30432 41497
rect 31576 41488 31628 41540
rect 31944 41599 31996 41608
rect 31944 41565 31953 41599
rect 31953 41565 31987 41599
rect 31987 41565 31996 41599
rect 31944 41556 31996 41565
rect 33876 41556 33928 41608
rect 36544 41599 36596 41608
rect 36544 41565 36553 41599
rect 36553 41565 36587 41599
rect 36587 41565 36596 41599
rect 36544 41556 36596 41565
rect 38384 41624 38436 41676
rect 43352 41692 43404 41744
rect 46388 41760 46440 41812
rect 47032 41803 47084 41812
rect 47032 41769 47041 41803
rect 47041 41769 47075 41803
rect 47075 41769 47084 41803
rect 47032 41760 47084 41769
rect 47216 41760 47268 41812
rect 49056 41803 49108 41812
rect 49056 41769 49065 41803
rect 49065 41769 49099 41803
rect 49099 41769 49108 41803
rect 49056 41760 49108 41769
rect 49516 41760 49568 41812
rect 50252 41803 50304 41812
rect 50252 41769 50261 41803
rect 50261 41769 50295 41803
rect 50295 41769 50304 41803
rect 50252 41760 50304 41769
rect 51540 41760 51592 41812
rect 51816 41760 51868 41812
rect 53472 41760 53524 41812
rect 45468 41692 45520 41744
rect 46020 41692 46072 41744
rect 46848 41692 46900 41744
rect 47492 41735 47544 41744
rect 47492 41701 47501 41735
rect 47501 41701 47535 41735
rect 47535 41701 47544 41735
rect 47492 41692 47544 41701
rect 47860 41692 47912 41744
rect 51448 41692 51500 41744
rect 52460 41735 52512 41744
rect 52460 41701 52469 41735
rect 52469 41701 52503 41735
rect 52503 41701 52512 41735
rect 52460 41692 52512 41701
rect 58348 41760 58400 41812
rect 41328 41624 41380 41676
rect 45100 41667 45152 41676
rect 45100 41633 45109 41667
rect 45109 41633 45143 41667
rect 45143 41633 45152 41667
rect 45100 41624 45152 41633
rect 37832 41556 37884 41608
rect 39856 41599 39908 41608
rect 39856 41565 39865 41599
rect 39865 41565 39899 41599
rect 39899 41565 39908 41599
rect 39856 41556 39908 41565
rect 40408 41556 40460 41608
rect 42708 41599 42760 41608
rect 42708 41565 42717 41599
rect 42717 41565 42751 41599
rect 42751 41565 42760 41599
rect 42708 41556 42760 41565
rect 42800 41556 42852 41608
rect 43352 41556 43404 41608
rect 44456 41556 44508 41608
rect 47952 41624 48004 41676
rect 48596 41624 48648 41676
rect 51356 41624 51408 41676
rect 55128 41624 55180 41676
rect 57704 41667 57756 41676
rect 57704 41633 57713 41667
rect 57713 41633 57747 41667
rect 57747 41633 57756 41667
rect 57704 41624 57756 41633
rect 31852 41488 31904 41540
rect 33508 41488 33560 41540
rect 34428 41488 34480 41540
rect 47584 41599 47636 41608
rect 47584 41565 47593 41599
rect 47593 41565 47627 41599
rect 47627 41565 47636 41599
rect 47584 41556 47636 41565
rect 48228 41488 48280 41540
rect 21732 41420 21784 41472
rect 23112 41420 23164 41472
rect 30472 41420 30524 41472
rect 30656 41420 30708 41472
rect 32036 41420 32088 41472
rect 32404 41420 32456 41472
rect 34520 41420 34572 41472
rect 34888 41463 34940 41472
rect 34888 41429 34897 41463
rect 34897 41429 34931 41463
rect 34931 41429 34940 41463
rect 34888 41420 34940 41429
rect 35900 41463 35952 41472
rect 35900 41429 35909 41463
rect 35909 41429 35943 41463
rect 35943 41429 35952 41463
rect 35900 41420 35952 41429
rect 37556 41463 37608 41472
rect 37556 41429 37565 41463
rect 37565 41429 37599 41463
rect 37599 41429 37608 41463
rect 37556 41420 37608 41429
rect 41696 41420 41748 41472
rect 47768 41420 47820 41472
rect 50804 41599 50856 41608
rect 50804 41565 50813 41599
rect 50813 41565 50847 41599
rect 50847 41565 50856 41599
rect 50804 41556 50856 41565
rect 49976 41488 50028 41540
rect 50896 41488 50948 41540
rect 56140 41599 56192 41608
rect 56140 41565 56149 41599
rect 56149 41565 56183 41599
rect 56183 41565 56192 41599
rect 56140 41556 56192 41565
rect 56508 41556 56560 41608
rect 54116 41488 54168 41540
rect 54944 41488 54996 41540
rect 55680 41420 55732 41472
rect 56416 41420 56468 41472
rect 57796 41420 57848 41472
rect 1998 41318 2050 41370
rect 2062 41318 2114 41370
rect 2126 41318 2178 41370
rect 2190 41318 2242 41370
rect 2254 41318 2306 41370
rect 50998 41318 51050 41370
rect 51062 41318 51114 41370
rect 51126 41318 51178 41370
rect 51190 41318 51242 41370
rect 51254 41318 51306 41370
rect 13728 41216 13780 41268
rect 15660 41216 15712 41268
rect 16764 41259 16816 41268
rect 16764 41225 16773 41259
rect 16773 41225 16807 41259
rect 16807 41225 16816 41259
rect 16764 41216 16816 41225
rect 20996 41216 21048 41268
rect 21548 41216 21600 41268
rect 23756 41216 23808 41268
rect 13084 41148 13136 41200
rect 8760 41080 8812 41132
rect 10048 41080 10100 41132
rect 11428 41123 11480 41132
rect 11428 41089 11437 41123
rect 11437 41089 11471 41123
rect 11471 41089 11480 41123
rect 11428 41080 11480 41089
rect 12440 41080 12492 41132
rect 14648 41148 14700 41200
rect 19156 41148 19208 41200
rect 21732 41191 21784 41200
rect 21732 41157 21741 41191
rect 21741 41157 21775 41191
rect 21775 41157 21784 41191
rect 21732 41148 21784 41157
rect 22560 41148 22612 41200
rect 13820 41012 13872 41064
rect 9680 40944 9732 40996
rect 9772 40944 9824 40996
rect 10140 40944 10192 40996
rect 11888 40987 11940 40996
rect 11888 40953 11897 40987
rect 11897 40953 11931 40987
rect 11931 40953 11940 40987
rect 11888 40944 11940 40953
rect 12900 40944 12952 40996
rect 17500 41123 17552 41132
rect 17500 41089 17509 41123
rect 17509 41089 17543 41123
rect 17543 41089 17552 41123
rect 17500 41080 17552 41089
rect 17868 41080 17920 41132
rect 17960 41080 18012 41132
rect 19984 41123 20036 41132
rect 19984 41089 19993 41123
rect 19993 41089 20027 41123
rect 20027 41089 20036 41123
rect 19984 41080 20036 41089
rect 20260 41123 20312 41132
rect 20260 41089 20269 41123
rect 20269 41089 20303 41123
rect 20303 41089 20312 41123
rect 20260 41080 20312 41089
rect 21456 41080 21508 41132
rect 25596 41216 25648 41268
rect 26240 41216 26292 41268
rect 26976 41216 27028 41268
rect 27160 41216 27212 41268
rect 25228 41148 25280 41200
rect 25872 41148 25924 41200
rect 33876 41259 33928 41268
rect 33876 41225 33885 41259
rect 33885 41225 33919 41259
rect 33919 41225 33928 41259
rect 33876 41216 33928 41225
rect 35808 41216 35860 41268
rect 37096 41216 37148 41268
rect 37832 41259 37884 41268
rect 37832 41225 37841 41259
rect 37841 41225 37875 41259
rect 37875 41225 37884 41259
rect 37832 41216 37884 41225
rect 39120 41216 39172 41268
rect 39488 41216 39540 41268
rect 24676 41123 24728 41132
rect 18052 41012 18104 41064
rect 19064 41012 19116 41064
rect 23020 41012 23072 41064
rect 24676 41089 24685 41123
rect 24685 41089 24719 41123
rect 24719 41089 24728 41123
rect 24676 41080 24728 41089
rect 25136 41080 25188 41132
rect 26884 41080 26936 41132
rect 31116 41080 31168 41132
rect 31576 41080 31628 41132
rect 24768 41012 24820 41064
rect 8944 40876 8996 40928
rect 11428 40876 11480 40928
rect 12808 40876 12860 40928
rect 15200 40944 15252 40996
rect 15292 40987 15344 40996
rect 15292 40953 15301 40987
rect 15301 40953 15335 40987
rect 15335 40953 15344 40987
rect 15292 40944 15344 40953
rect 16304 40944 16356 40996
rect 18788 40944 18840 40996
rect 13820 40919 13872 40928
rect 13820 40885 13829 40919
rect 13829 40885 13863 40919
rect 13863 40885 13872 40919
rect 13820 40876 13872 40885
rect 14096 40876 14148 40928
rect 14464 40876 14516 40928
rect 16948 40876 17000 40928
rect 17408 40876 17460 40928
rect 20352 40944 20404 40996
rect 27068 41055 27120 41064
rect 27068 41021 27077 41055
rect 27077 41021 27111 41055
rect 27111 41021 27120 41055
rect 27068 41012 27120 41021
rect 27436 41012 27488 41064
rect 30104 41012 30156 41064
rect 30656 41055 30708 41064
rect 30656 41021 30665 41055
rect 30665 41021 30699 41055
rect 30699 41021 30708 41055
rect 30656 41012 30708 41021
rect 32128 41123 32180 41132
rect 32128 41089 32137 41123
rect 32137 41089 32171 41123
rect 32171 41089 32180 41123
rect 32128 41080 32180 41089
rect 34244 41080 34296 41132
rect 35256 41080 35308 41132
rect 35716 41080 35768 41132
rect 35900 41080 35952 41132
rect 31852 40944 31904 40996
rect 34888 41012 34940 41064
rect 47860 41259 47912 41268
rect 47860 41225 47869 41259
rect 47869 41225 47903 41259
rect 47903 41225 47912 41259
rect 47860 41216 47912 41225
rect 48596 41259 48648 41268
rect 48596 41225 48605 41259
rect 48605 41225 48639 41259
rect 48639 41225 48648 41259
rect 48596 41216 48648 41225
rect 52276 41216 52328 41268
rect 38936 41148 38988 41200
rect 39764 41123 39816 41132
rect 39764 41089 39773 41123
rect 39773 41089 39807 41123
rect 39807 41089 39816 41123
rect 39764 41080 39816 41089
rect 40132 41148 40184 41200
rect 40684 41148 40736 41200
rect 42708 41148 42760 41200
rect 22192 40919 22244 40928
rect 22192 40885 22201 40919
rect 22201 40885 22235 40919
rect 22235 40885 22244 40919
rect 22192 40876 22244 40885
rect 22284 40919 22336 40928
rect 22284 40885 22293 40919
rect 22293 40885 22327 40919
rect 22327 40885 22336 40919
rect 22284 40876 22336 40885
rect 24400 40876 24452 40928
rect 24676 40876 24728 40928
rect 24860 40876 24912 40928
rect 27528 40876 27580 40928
rect 29092 40876 29144 40928
rect 29920 40876 29972 40928
rect 32220 40876 32272 40928
rect 34152 40944 34204 40996
rect 35900 40987 35952 40996
rect 35900 40953 35909 40987
rect 35909 40953 35943 40987
rect 35943 40953 35952 40987
rect 35900 40944 35952 40953
rect 36268 40944 36320 40996
rect 33416 40876 33468 40928
rect 34612 40919 34664 40928
rect 34612 40885 34621 40919
rect 34621 40885 34655 40919
rect 34655 40885 34664 40919
rect 34612 40876 34664 40885
rect 35072 40876 35124 40928
rect 35440 40919 35492 40928
rect 35440 40885 35449 40919
rect 35449 40885 35483 40919
rect 35483 40885 35492 40919
rect 35440 40876 35492 40885
rect 37188 41012 37240 41064
rect 37096 40944 37148 40996
rect 43076 41080 43128 41132
rect 46112 41148 46164 41200
rect 52552 41148 52604 41200
rect 53196 41216 53248 41268
rect 57704 41216 57756 41268
rect 41972 41055 42024 41064
rect 41972 41021 41981 41055
rect 41981 41021 42015 41055
rect 42015 41021 42024 41055
rect 41972 41012 42024 41021
rect 42800 41012 42852 41064
rect 45008 41012 45060 41064
rect 47860 41080 47912 41132
rect 47952 41123 48004 41132
rect 47952 41089 47961 41123
rect 47961 41089 47995 41123
rect 47995 41089 48004 41123
rect 47952 41080 48004 41089
rect 48780 41080 48832 41132
rect 49332 41080 49384 41132
rect 50620 41080 50672 41132
rect 54024 41148 54076 41200
rect 53656 41123 53708 41132
rect 53656 41089 53665 41123
rect 53665 41089 53699 41123
rect 53699 41089 53708 41123
rect 53656 41080 53708 41089
rect 54484 41148 54536 41200
rect 54852 41148 54904 41200
rect 54208 41080 54260 41132
rect 55036 41080 55088 41132
rect 41420 40944 41472 40996
rect 41604 40944 41656 40996
rect 41696 40987 41748 40996
rect 41696 40953 41705 40987
rect 41705 40953 41739 40987
rect 41739 40953 41748 40987
rect 41696 40944 41748 40953
rect 42248 40944 42300 40996
rect 43168 40944 43220 40996
rect 45100 40944 45152 40996
rect 45468 40944 45520 40996
rect 40040 40876 40092 40928
rect 40408 40876 40460 40928
rect 40960 40876 41012 40928
rect 42800 40876 42852 40928
rect 42892 40919 42944 40928
rect 42892 40885 42901 40919
rect 42901 40885 42935 40919
rect 42935 40885 42944 40919
rect 42892 40876 42944 40885
rect 43076 40876 43128 40928
rect 46112 40876 46164 40928
rect 46480 40944 46532 40996
rect 47492 40987 47544 40996
rect 47492 40953 47501 40987
rect 47501 40953 47535 40987
rect 47535 40953 47544 40987
rect 47492 40944 47544 40953
rect 48044 40944 48096 40996
rect 49516 40944 49568 40996
rect 49608 40944 49660 40996
rect 51080 41012 51132 41064
rect 51172 41055 51224 41064
rect 51172 41021 51181 41055
rect 51181 41021 51215 41055
rect 51215 41021 51224 41055
rect 51172 41012 51224 41021
rect 56416 41012 56468 41064
rect 56692 41123 56744 41132
rect 56692 41089 56701 41123
rect 56701 41089 56735 41123
rect 56735 41089 56744 41123
rect 56692 41080 56744 41089
rect 57060 41080 57112 41132
rect 46296 40919 46348 40928
rect 46296 40885 46305 40919
rect 46305 40885 46339 40919
rect 46339 40885 46348 40919
rect 46296 40876 46348 40885
rect 46664 40919 46716 40928
rect 46664 40885 46673 40919
rect 46673 40885 46707 40919
rect 46707 40885 46716 40919
rect 46664 40876 46716 40885
rect 49424 40876 49476 40928
rect 50160 40919 50212 40928
rect 50160 40885 50169 40919
rect 50169 40885 50203 40919
rect 50203 40885 50212 40919
rect 50160 40876 50212 40885
rect 51356 40876 51408 40928
rect 52368 40876 52420 40928
rect 52828 40876 52880 40928
rect 54760 40944 54812 40996
rect 55036 40876 55088 40928
rect 55220 40876 55272 40928
rect 55680 40919 55732 40928
rect 55680 40885 55689 40919
rect 55689 40885 55723 40919
rect 55723 40885 55732 40919
rect 55680 40876 55732 40885
rect 55772 40919 55824 40928
rect 55772 40885 55781 40919
rect 55781 40885 55815 40919
rect 55815 40885 55824 40919
rect 55772 40876 55824 40885
rect 56140 40919 56192 40928
rect 56140 40885 56149 40919
rect 56149 40885 56183 40919
rect 56183 40885 56192 40919
rect 56140 40876 56192 40885
rect 56600 40987 56652 40996
rect 56600 40953 56609 40987
rect 56609 40953 56643 40987
rect 56643 40953 56652 40987
rect 56600 40944 56652 40953
rect 57060 40987 57112 40996
rect 57060 40953 57069 40987
rect 57069 40953 57103 40987
rect 57103 40953 57112 40987
rect 57060 40944 57112 40953
rect 57152 40919 57204 40928
rect 57152 40885 57161 40919
rect 57161 40885 57195 40919
rect 57195 40885 57204 40919
rect 57152 40876 57204 40885
rect 57612 41055 57664 41064
rect 57612 41021 57621 41055
rect 57621 41021 57655 41055
rect 57655 41021 57664 41055
rect 57612 41012 57664 41021
rect 57520 40944 57572 40996
rect 66076 41012 66128 41064
rect 64880 40876 64932 40928
rect 2918 40774 2970 40826
rect 2982 40774 3034 40826
rect 3046 40774 3098 40826
rect 3110 40774 3162 40826
rect 3174 40774 3226 40826
rect 51918 40774 51970 40826
rect 51982 40774 52034 40826
rect 52046 40774 52098 40826
rect 52110 40774 52162 40826
rect 52174 40774 52226 40826
rect 10692 40672 10744 40724
rect 11428 40672 11480 40724
rect 16948 40672 17000 40724
rect 10140 40536 10192 40588
rect 10324 40536 10376 40588
rect 11428 40579 11480 40588
rect 11428 40545 11437 40579
rect 11437 40545 11471 40579
rect 11471 40545 11480 40579
rect 11428 40536 11480 40545
rect 8760 40511 8812 40520
rect 8760 40477 8769 40511
rect 8769 40477 8803 40511
rect 8803 40477 8812 40511
rect 8760 40468 8812 40477
rect 9036 40511 9088 40520
rect 9036 40477 9045 40511
rect 9045 40477 9079 40511
rect 9079 40477 9088 40511
rect 9036 40468 9088 40477
rect 9772 40468 9824 40520
rect 14096 40647 14148 40656
rect 14096 40613 14105 40647
rect 14105 40613 14139 40647
rect 14139 40613 14148 40647
rect 14096 40604 14148 40613
rect 15200 40536 15252 40588
rect 12256 40468 12308 40520
rect 13728 40468 13780 40520
rect 15384 40511 15436 40520
rect 15384 40477 15393 40511
rect 15393 40477 15427 40511
rect 15427 40477 15436 40511
rect 15384 40468 15436 40477
rect 16764 40604 16816 40656
rect 17408 40604 17460 40656
rect 17960 40536 18012 40588
rect 20812 40672 20864 40724
rect 21272 40715 21324 40724
rect 21272 40681 21281 40715
rect 21281 40681 21315 40715
rect 21315 40681 21324 40715
rect 21272 40672 21324 40681
rect 22192 40715 22244 40724
rect 22192 40681 22201 40715
rect 22201 40681 22235 40715
rect 22235 40681 22244 40715
rect 22192 40672 22244 40681
rect 24768 40672 24820 40724
rect 26240 40672 26292 40724
rect 23940 40647 23992 40656
rect 23940 40613 23949 40647
rect 23949 40613 23983 40647
rect 23983 40613 23992 40647
rect 23940 40604 23992 40613
rect 25228 40604 25280 40656
rect 16764 40468 16816 40520
rect 17500 40468 17552 40520
rect 18052 40468 18104 40520
rect 20444 40536 20496 40588
rect 22836 40579 22888 40588
rect 22836 40545 22845 40579
rect 22845 40545 22879 40579
rect 22879 40545 22888 40579
rect 22836 40536 22888 40545
rect 26424 40536 26476 40588
rect 26516 40536 26568 40588
rect 29092 40715 29144 40724
rect 29092 40681 29101 40715
rect 29101 40681 29135 40715
rect 29135 40681 29144 40715
rect 29092 40672 29144 40681
rect 29920 40647 29972 40656
rect 29920 40613 29929 40647
rect 29929 40613 29963 40647
rect 29963 40613 29972 40647
rect 29920 40604 29972 40613
rect 30012 40604 30064 40656
rect 30564 40672 30616 40724
rect 30656 40672 30708 40724
rect 33232 40672 33284 40724
rect 33692 40672 33744 40724
rect 34612 40672 34664 40724
rect 32128 40604 32180 40656
rect 33048 40604 33100 40656
rect 35900 40672 35952 40724
rect 36544 40715 36596 40724
rect 36544 40681 36553 40715
rect 36553 40681 36587 40715
rect 36587 40681 36596 40715
rect 36544 40672 36596 40681
rect 38568 40672 38620 40724
rect 28816 40536 28868 40588
rect 31668 40579 31720 40588
rect 31668 40545 31677 40579
rect 31677 40545 31711 40579
rect 31711 40545 31720 40579
rect 31668 40536 31720 40545
rect 33140 40536 33192 40588
rect 18328 40511 18380 40520
rect 18328 40477 18337 40511
rect 18337 40477 18371 40511
rect 18371 40477 18380 40511
rect 18328 40468 18380 40477
rect 18420 40511 18472 40520
rect 18420 40477 18429 40511
rect 18429 40477 18463 40511
rect 18463 40477 18472 40511
rect 18420 40468 18472 40477
rect 19340 40511 19392 40520
rect 19340 40477 19349 40511
rect 19349 40477 19383 40511
rect 19383 40477 19392 40511
rect 19340 40468 19392 40477
rect 19892 40468 19944 40520
rect 20352 40468 20404 40520
rect 20720 40468 20772 40520
rect 21456 40468 21508 40520
rect 15568 40332 15620 40384
rect 16856 40375 16908 40384
rect 16856 40341 16865 40375
rect 16865 40341 16899 40375
rect 16899 40341 16908 40375
rect 16856 40332 16908 40341
rect 17776 40332 17828 40384
rect 21640 40400 21692 40452
rect 20628 40332 20680 40384
rect 22192 40468 22244 40520
rect 23572 40511 23624 40520
rect 23572 40477 23581 40511
rect 23581 40477 23615 40511
rect 23615 40477 23624 40511
rect 23572 40468 23624 40477
rect 23664 40511 23716 40520
rect 23664 40477 23673 40511
rect 23673 40477 23707 40511
rect 23707 40477 23716 40511
rect 23664 40468 23716 40477
rect 25136 40468 25188 40520
rect 22100 40332 22152 40384
rect 22928 40375 22980 40384
rect 22928 40341 22937 40375
rect 22937 40341 22971 40375
rect 22971 40341 22980 40375
rect 22928 40332 22980 40341
rect 23296 40332 23348 40384
rect 26332 40468 26384 40520
rect 26792 40468 26844 40520
rect 26884 40511 26936 40520
rect 26884 40477 26893 40511
rect 26893 40477 26927 40511
rect 26927 40477 26936 40511
rect 26884 40468 26936 40477
rect 27068 40511 27120 40520
rect 27068 40477 27077 40511
rect 27077 40477 27111 40511
rect 27111 40477 27120 40511
rect 27068 40468 27120 40477
rect 27528 40468 27580 40520
rect 29276 40468 29328 40520
rect 29368 40468 29420 40520
rect 30380 40468 30432 40520
rect 26148 40400 26200 40452
rect 31208 40468 31260 40520
rect 31852 40468 31904 40520
rect 32956 40468 33008 40520
rect 33784 40536 33836 40588
rect 35072 40647 35124 40656
rect 35072 40613 35081 40647
rect 35081 40613 35115 40647
rect 35115 40613 35124 40647
rect 35072 40604 35124 40613
rect 35532 40604 35584 40656
rect 37556 40604 37608 40656
rect 39028 40604 39080 40656
rect 37188 40536 37240 40588
rect 40040 40604 40092 40656
rect 40776 40604 40828 40656
rect 41328 40604 41380 40656
rect 51172 40672 51224 40724
rect 51448 40672 51500 40724
rect 52368 40672 52420 40724
rect 44732 40604 44784 40656
rect 33508 40468 33560 40520
rect 33968 40511 34020 40520
rect 33968 40477 33977 40511
rect 33977 40477 34011 40511
rect 34011 40477 34020 40511
rect 33968 40468 34020 40477
rect 34060 40511 34112 40520
rect 34060 40477 34069 40511
rect 34069 40477 34103 40511
rect 34103 40477 34112 40511
rect 34060 40468 34112 40477
rect 36084 40468 36136 40520
rect 37648 40468 37700 40520
rect 38384 40468 38436 40520
rect 40132 40536 40184 40588
rect 40960 40536 41012 40588
rect 39304 40468 39356 40520
rect 39856 40468 39908 40520
rect 25596 40332 25648 40384
rect 26700 40332 26752 40384
rect 28080 40375 28132 40384
rect 28080 40341 28089 40375
rect 28089 40341 28123 40375
rect 28123 40341 28132 40375
rect 28080 40332 28132 40341
rect 29276 40332 29328 40384
rect 30472 40332 30524 40384
rect 31852 40332 31904 40384
rect 32128 40375 32180 40384
rect 32128 40341 32137 40375
rect 32137 40341 32171 40375
rect 32171 40341 32180 40375
rect 32128 40332 32180 40341
rect 40316 40443 40368 40452
rect 40316 40409 40325 40443
rect 40325 40409 40359 40443
rect 40359 40409 40368 40443
rect 40316 40400 40368 40409
rect 40684 40400 40736 40452
rect 38660 40332 38712 40384
rect 39212 40375 39264 40384
rect 39212 40341 39221 40375
rect 39221 40341 39255 40375
rect 39255 40341 39264 40375
rect 39212 40332 39264 40341
rect 40408 40332 40460 40384
rect 41972 40536 42024 40588
rect 45468 40579 45520 40588
rect 45468 40545 45477 40579
rect 45477 40545 45511 40579
rect 45511 40545 45520 40579
rect 45468 40536 45520 40545
rect 45744 40604 45796 40656
rect 46388 40604 46440 40656
rect 49424 40647 49476 40656
rect 49424 40613 49433 40647
rect 49433 40613 49467 40647
rect 49467 40613 49476 40647
rect 49424 40604 49476 40613
rect 49976 40604 50028 40656
rect 50712 40604 50764 40656
rect 46204 40536 46256 40588
rect 47676 40536 47728 40588
rect 47768 40536 47820 40588
rect 48228 40536 48280 40588
rect 51080 40536 51132 40588
rect 52276 40536 52328 40588
rect 43720 40511 43772 40520
rect 43720 40477 43729 40511
rect 43729 40477 43763 40511
rect 43763 40477 43772 40511
rect 43720 40468 43772 40477
rect 43352 40375 43404 40384
rect 43352 40341 43361 40375
rect 43361 40341 43395 40375
rect 43395 40341 43404 40375
rect 43352 40332 43404 40341
rect 47860 40468 47912 40520
rect 48504 40511 48556 40520
rect 48504 40477 48513 40511
rect 48513 40477 48547 40511
rect 48547 40477 48556 40511
rect 48504 40468 48556 40477
rect 47400 40400 47452 40452
rect 48228 40400 48280 40452
rect 50160 40468 50212 40520
rect 50712 40468 50764 40520
rect 51816 40511 51868 40520
rect 51816 40477 51825 40511
rect 51825 40477 51859 40511
rect 51859 40477 51868 40511
rect 51816 40468 51868 40477
rect 52828 40511 52880 40520
rect 52828 40477 52837 40511
rect 52837 40477 52871 40511
rect 52871 40477 52880 40511
rect 52828 40468 52880 40477
rect 53472 40536 53524 40588
rect 55128 40672 55180 40724
rect 55220 40647 55272 40656
rect 55220 40613 55229 40647
rect 55229 40613 55263 40647
rect 55263 40613 55272 40647
rect 55220 40604 55272 40613
rect 56692 40672 56744 40724
rect 57520 40672 57572 40724
rect 57704 40672 57756 40724
rect 60648 40672 60700 40724
rect 54208 40468 54260 40520
rect 54576 40511 54628 40520
rect 54576 40477 54585 40511
rect 54585 40477 54619 40511
rect 54619 40477 54628 40511
rect 54576 40468 54628 40477
rect 55772 40468 55824 40520
rect 47768 40332 47820 40384
rect 49056 40375 49108 40384
rect 49056 40341 49065 40375
rect 49065 40341 49099 40375
rect 49099 40341 49108 40375
rect 49056 40332 49108 40341
rect 51356 40400 51408 40452
rect 53564 40332 53616 40384
rect 54484 40332 54536 40384
rect 56692 40332 56744 40384
rect 1998 40230 2050 40282
rect 2062 40230 2114 40282
rect 2126 40230 2178 40282
rect 2190 40230 2242 40282
rect 2254 40230 2306 40282
rect 50998 40230 51050 40282
rect 51062 40230 51114 40282
rect 51126 40230 51178 40282
rect 51190 40230 51242 40282
rect 51254 40230 51306 40282
rect 9036 40128 9088 40180
rect 9312 40035 9364 40044
rect 9312 40001 9321 40035
rect 9321 40001 9355 40035
rect 9355 40001 9364 40035
rect 9312 39992 9364 40001
rect 10324 40060 10376 40112
rect 10416 39992 10468 40044
rect 10968 40128 11020 40180
rect 12808 39992 12860 40044
rect 14188 40035 14240 40044
rect 14188 40001 14197 40035
rect 14197 40001 14231 40035
rect 14231 40001 14240 40035
rect 14188 39992 14240 40001
rect 14464 40035 14516 40044
rect 14464 40001 14473 40035
rect 14473 40001 14507 40035
rect 14507 40001 14516 40035
rect 14464 39992 14516 40001
rect 15200 39992 15252 40044
rect 16856 40128 16908 40180
rect 19800 40128 19852 40180
rect 20444 40128 20496 40180
rect 22284 40128 22336 40180
rect 23940 40128 23992 40180
rect 21088 40060 21140 40112
rect 17316 39992 17368 40044
rect 17960 39992 18012 40044
rect 20076 39992 20128 40044
rect 21640 40060 21692 40112
rect 22192 40060 22244 40112
rect 22100 39992 22152 40044
rect 22560 40035 22612 40044
rect 22560 40001 22569 40035
rect 22569 40001 22603 40035
rect 22603 40001 22612 40035
rect 22560 39992 22612 40001
rect 23296 40060 23348 40112
rect 24492 40060 24544 40112
rect 26516 40128 26568 40180
rect 26700 40171 26752 40180
rect 26700 40137 26721 40171
rect 26721 40137 26752 40171
rect 26700 40128 26752 40137
rect 24400 39992 24452 40044
rect 27988 40128 28040 40180
rect 28816 40171 28868 40180
rect 28816 40137 28825 40171
rect 28825 40137 28859 40171
rect 28859 40137 28868 40171
rect 28816 40128 28868 40137
rect 26976 40060 27028 40112
rect 30288 40128 30340 40180
rect 30472 40128 30524 40180
rect 36084 40128 36136 40180
rect 36268 40128 36320 40180
rect 36728 40128 36780 40180
rect 7932 39924 7984 39976
rect 12440 39924 12492 39976
rect 13728 39924 13780 39976
rect 20996 39924 21048 39976
rect 22928 39924 22980 39976
rect 23572 39924 23624 39976
rect 24216 39924 24268 39976
rect 25412 39924 25464 39976
rect 29368 39992 29420 40044
rect 31576 40060 31628 40112
rect 35256 40060 35308 40112
rect 39212 40128 39264 40180
rect 39396 40128 39448 40180
rect 41604 40128 41656 40180
rect 41880 40128 41932 40180
rect 46296 40128 46348 40180
rect 30104 39992 30156 40044
rect 30564 39992 30616 40044
rect 31300 39992 31352 40044
rect 31392 39992 31444 40044
rect 36452 39992 36504 40044
rect 37188 39992 37240 40044
rect 38292 39992 38344 40044
rect 8944 39856 8996 39908
rect 8208 39788 8260 39840
rect 9680 39788 9732 39840
rect 10140 39788 10192 39840
rect 10692 39831 10744 39840
rect 10692 39797 10701 39831
rect 10701 39797 10735 39831
rect 10735 39797 10744 39831
rect 10692 39788 10744 39797
rect 11060 39788 11112 39840
rect 11428 39856 11480 39908
rect 16304 39856 16356 39908
rect 11612 39831 11664 39840
rect 11612 39797 11621 39831
rect 11621 39797 11655 39831
rect 11655 39797 11664 39831
rect 11612 39788 11664 39797
rect 12624 39831 12676 39840
rect 12624 39797 12633 39831
rect 12633 39797 12667 39831
rect 12667 39797 12676 39831
rect 12624 39788 12676 39797
rect 18328 39856 18380 39908
rect 19892 39856 19944 39908
rect 18052 39788 18104 39840
rect 18512 39788 18564 39840
rect 19064 39831 19116 39840
rect 19064 39797 19073 39831
rect 19073 39797 19107 39831
rect 19107 39797 19116 39831
rect 19064 39788 19116 39797
rect 19156 39788 19208 39840
rect 24952 39856 25004 39908
rect 22744 39788 22796 39840
rect 24676 39788 24728 39840
rect 26056 39788 26108 39840
rect 39028 39924 39080 39976
rect 39488 40035 39540 40044
rect 39488 40001 39497 40035
rect 39497 40001 39531 40035
rect 39531 40001 39540 40035
rect 39488 39992 39540 40001
rect 40132 40035 40184 40044
rect 40132 40001 40141 40035
rect 40141 40001 40175 40035
rect 40175 40001 40184 40035
rect 40132 39992 40184 40001
rect 40224 39992 40276 40044
rect 43076 39992 43128 40044
rect 43720 39992 43772 40044
rect 44088 39992 44140 40044
rect 48044 40128 48096 40180
rect 48504 40128 48556 40180
rect 49608 40171 49660 40180
rect 49608 40137 49617 40171
rect 49617 40137 49651 40171
rect 49651 40137 49660 40171
rect 49608 40128 49660 40137
rect 47768 40060 47820 40112
rect 47400 39992 47452 40044
rect 49516 40060 49568 40112
rect 51816 40128 51868 40180
rect 56600 40128 56652 40180
rect 57520 40128 57572 40180
rect 57152 40060 57204 40112
rect 40868 39967 40920 39976
rect 40868 39933 40877 39967
rect 40877 39933 40911 39967
rect 40911 39933 40920 39967
rect 40868 39924 40920 39933
rect 42432 39924 42484 39976
rect 45376 39924 45428 39976
rect 27344 39899 27396 39908
rect 27344 39865 27353 39899
rect 27353 39865 27387 39899
rect 27387 39865 27396 39899
rect 27344 39856 27396 39865
rect 28632 39856 28684 39908
rect 29828 39856 29880 39908
rect 30380 39856 30432 39908
rect 30564 39856 30616 39908
rect 32588 39856 32640 39908
rect 33324 39856 33376 39908
rect 35532 39856 35584 39908
rect 36820 39899 36872 39908
rect 36820 39865 36829 39899
rect 36829 39865 36863 39899
rect 36863 39865 36872 39899
rect 36820 39856 36872 39865
rect 27436 39788 27488 39840
rect 28908 39788 28960 39840
rect 30748 39788 30800 39840
rect 31576 39831 31628 39840
rect 31576 39797 31585 39831
rect 31585 39797 31619 39831
rect 31619 39797 31628 39831
rect 31576 39788 31628 39797
rect 32956 39831 33008 39840
rect 32956 39797 32965 39831
rect 32965 39797 32999 39831
rect 32999 39797 33008 39831
rect 32956 39788 33008 39797
rect 35256 39788 35308 39840
rect 35992 39788 36044 39840
rect 37280 39788 37332 39840
rect 39028 39788 39080 39840
rect 39396 39788 39448 39840
rect 39672 39788 39724 39840
rect 39856 39788 39908 39840
rect 41420 39856 41472 39908
rect 41880 39856 41932 39908
rect 46204 39856 46256 39908
rect 42892 39788 42944 39840
rect 43260 39788 43312 39840
rect 43536 39831 43588 39840
rect 43536 39797 43545 39831
rect 43545 39797 43579 39831
rect 43579 39797 43588 39831
rect 43536 39788 43588 39797
rect 45192 39831 45244 39840
rect 45192 39797 45201 39831
rect 45201 39797 45235 39831
rect 45235 39797 45244 39831
rect 45192 39788 45244 39797
rect 46480 39788 46532 39840
rect 46664 39856 46716 39908
rect 48412 39924 48464 39976
rect 49056 39967 49108 39976
rect 49056 39933 49065 39967
rect 49065 39933 49099 39967
rect 49099 39933 49108 39967
rect 49056 39924 49108 39933
rect 52460 39992 52512 40044
rect 53656 39992 53708 40044
rect 55680 40035 55732 40044
rect 55680 40001 55689 40035
rect 55689 40001 55723 40035
rect 55723 40001 55732 40035
rect 55680 39992 55732 40001
rect 58716 40060 58768 40112
rect 49976 39924 50028 39976
rect 47400 39788 47452 39840
rect 48596 39831 48648 39840
rect 48596 39797 48605 39831
rect 48605 39797 48639 39831
rect 48639 39797 48648 39831
rect 48596 39788 48648 39797
rect 48964 39831 49016 39840
rect 48964 39797 48973 39831
rect 48973 39797 49007 39831
rect 49007 39797 49016 39831
rect 48964 39788 49016 39797
rect 49792 39856 49844 39908
rect 50160 39788 50212 39840
rect 50896 39788 50948 39840
rect 53748 39924 53800 39976
rect 57704 39967 57756 39976
rect 57704 39933 57713 39967
rect 57713 39933 57747 39967
rect 57747 39933 57756 39967
rect 57704 39924 57756 39933
rect 52828 39856 52880 39908
rect 55312 39856 55364 39908
rect 57336 39856 57388 39908
rect 58808 39856 58860 39908
rect 55220 39788 55272 39840
rect 55772 39788 55824 39840
rect 57244 39831 57296 39840
rect 57244 39797 57253 39831
rect 57253 39797 57287 39831
rect 57287 39797 57296 39831
rect 57244 39788 57296 39797
rect 58072 39831 58124 39840
rect 58072 39797 58081 39831
rect 58081 39797 58115 39831
rect 58115 39797 58124 39831
rect 58072 39788 58124 39797
rect 58440 39831 58492 39840
rect 58440 39797 58449 39831
rect 58449 39797 58483 39831
rect 58483 39797 58492 39831
rect 58440 39788 58492 39797
rect 58900 39788 58952 39840
rect 2918 39686 2970 39738
rect 2982 39686 3034 39738
rect 3046 39686 3098 39738
rect 3110 39686 3162 39738
rect 3174 39686 3226 39738
rect 51918 39686 51970 39738
rect 51982 39686 52034 39738
rect 52046 39686 52098 39738
rect 52110 39686 52162 39738
rect 52174 39686 52226 39738
rect 9680 39516 9732 39568
rect 10140 39559 10192 39568
rect 10140 39525 10149 39559
rect 10149 39525 10183 39559
rect 10183 39525 10192 39559
rect 10140 39516 10192 39525
rect 14188 39584 14240 39636
rect 15292 39584 15344 39636
rect 15568 39627 15620 39636
rect 15568 39593 15577 39627
rect 15577 39593 15611 39627
rect 15611 39593 15620 39627
rect 15568 39584 15620 39593
rect 16488 39584 16540 39636
rect 17960 39584 18012 39636
rect 19156 39584 19208 39636
rect 20076 39627 20128 39636
rect 20076 39593 20085 39627
rect 20085 39593 20119 39627
rect 20119 39593 20128 39627
rect 20076 39584 20128 39593
rect 21548 39584 21600 39636
rect 12900 39516 12952 39568
rect 14556 39516 14608 39568
rect 17776 39516 17828 39568
rect 18788 39559 18840 39568
rect 18788 39525 18797 39559
rect 18797 39525 18831 39559
rect 18831 39525 18840 39559
rect 18788 39516 18840 39525
rect 19064 39516 19116 39568
rect 11336 39491 11388 39500
rect 11336 39457 11345 39491
rect 11345 39457 11379 39491
rect 11379 39457 11388 39491
rect 11336 39448 11388 39457
rect 12072 39448 12124 39500
rect 15108 39448 15160 39500
rect 17500 39491 17552 39500
rect 17500 39457 17509 39491
rect 17509 39457 17543 39491
rect 17543 39457 17552 39491
rect 17500 39448 17552 39457
rect 18052 39448 18104 39500
rect 20628 39448 20680 39500
rect 21640 39491 21692 39500
rect 21640 39457 21649 39491
rect 21649 39457 21683 39491
rect 21683 39457 21692 39491
rect 21640 39448 21692 39457
rect 22744 39559 22796 39568
rect 22744 39525 22753 39559
rect 22753 39525 22787 39559
rect 22787 39525 22796 39559
rect 22744 39516 22796 39525
rect 25044 39584 25096 39636
rect 25596 39584 25648 39636
rect 26148 39584 26200 39636
rect 26240 39627 26292 39636
rect 26240 39593 26249 39627
rect 26249 39593 26283 39627
rect 26283 39593 26292 39627
rect 26240 39584 26292 39593
rect 26424 39627 26476 39636
rect 26424 39593 26433 39627
rect 26433 39593 26467 39627
rect 26467 39593 26476 39627
rect 26424 39584 26476 39593
rect 26516 39584 26568 39636
rect 26976 39584 27028 39636
rect 27344 39584 27396 39636
rect 28080 39627 28132 39636
rect 28080 39593 28089 39627
rect 28089 39593 28123 39627
rect 28123 39593 28132 39627
rect 28080 39584 28132 39593
rect 24768 39559 24820 39568
rect 24768 39525 24777 39559
rect 24777 39525 24811 39559
rect 24811 39525 24820 39559
rect 24768 39516 24820 39525
rect 26056 39516 26108 39568
rect 27620 39516 27672 39568
rect 8208 39380 8260 39432
rect 11612 39423 11664 39432
rect 11612 39389 11621 39423
rect 11621 39389 11655 39423
rect 11655 39389 11664 39423
rect 11612 39380 11664 39389
rect 10416 39312 10468 39364
rect 7840 39287 7892 39296
rect 7840 39253 7849 39287
rect 7849 39253 7883 39287
rect 7883 39253 7892 39287
rect 7840 39244 7892 39253
rect 10324 39244 10376 39296
rect 12532 39380 12584 39432
rect 13820 39312 13872 39364
rect 16764 39380 16816 39432
rect 17316 39380 17368 39432
rect 15384 39312 15436 39364
rect 12440 39244 12492 39296
rect 13544 39244 13596 39296
rect 13912 39287 13964 39296
rect 13912 39253 13921 39287
rect 13921 39253 13955 39287
rect 13955 39253 13964 39287
rect 13912 39244 13964 39253
rect 14004 39287 14056 39296
rect 14004 39253 14013 39287
rect 14013 39253 14047 39287
rect 14047 39253 14056 39287
rect 14004 39244 14056 39253
rect 16856 39244 16908 39296
rect 18880 39380 18932 39432
rect 21364 39380 21416 39432
rect 21824 39423 21876 39432
rect 21824 39389 21833 39423
rect 21833 39389 21867 39423
rect 21867 39389 21876 39423
rect 21824 39380 21876 39389
rect 24216 39423 24268 39432
rect 24216 39389 24225 39423
rect 24225 39389 24259 39423
rect 24259 39389 24268 39423
rect 24216 39380 24268 39389
rect 25228 39380 25280 39432
rect 26240 39448 26292 39500
rect 26148 39380 26200 39432
rect 26516 39380 26568 39432
rect 27252 39448 27304 39500
rect 27436 39491 27488 39500
rect 27436 39457 27445 39491
rect 27445 39457 27479 39491
rect 27479 39457 27488 39491
rect 27436 39448 27488 39457
rect 28172 39423 28224 39432
rect 28172 39389 28181 39423
rect 28181 39389 28215 39423
rect 28215 39389 28224 39423
rect 28172 39380 28224 39389
rect 18420 39312 18472 39364
rect 19984 39312 20036 39364
rect 20628 39312 20680 39364
rect 20812 39312 20864 39364
rect 19892 39244 19944 39296
rect 26792 39312 26844 39364
rect 29736 39584 29788 39636
rect 30380 39627 30432 39636
rect 30380 39593 30389 39627
rect 30389 39593 30423 39627
rect 30423 39593 30432 39627
rect 30380 39584 30432 39593
rect 31300 39584 31352 39636
rect 32588 39584 32640 39636
rect 33140 39584 33192 39636
rect 33968 39584 34020 39636
rect 28908 39516 28960 39568
rect 30104 39516 30156 39568
rect 32128 39516 32180 39568
rect 29920 39448 29972 39500
rect 28816 39380 28868 39432
rect 30472 39448 30524 39500
rect 31944 39491 31996 39500
rect 31944 39457 31953 39491
rect 31953 39457 31987 39491
rect 31987 39457 31996 39491
rect 31944 39448 31996 39457
rect 34336 39491 34388 39500
rect 34336 39457 34345 39491
rect 34345 39457 34379 39491
rect 34379 39457 34388 39491
rect 34336 39448 34388 39457
rect 35440 39584 35492 39636
rect 36820 39584 36872 39636
rect 36912 39584 36964 39636
rect 39672 39584 39724 39636
rect 40040 39584 40092 39636
rect 40776 39584 40828 39636
rect 40960 39584 41012 39636
rect 42248 39627 42300 39636
rect 42248 39593 42257 39627
rect 42257 39593 42291 39627
rect 42291 39593 42300 39627
rect 42248 39584 42300 39593
rect 43076 39584 43128 39636
rect 35072 39516 35124 39568
rect 36544 39516 36596 39568
rect 39396 39516 39448 39568
rect 39856 39559 39908 39568
rect 39856 39525 39865 39559
rect 39865 39525 39899 39559
rect 39899 39525 39908 39559
rect 39856 39516 39908 39525
rect 43444 39516 43496 39568
rect 43812 39516 43864 39568
rect 30380 39312 30432 39364
rect 30840 39423 30892 39432
rect 30840 39389 30849 39423
rect 30849 39389 30883 39423
rect 30883 39389 30892 39423
rect 30840 39380 30892 39389
rect 31208 39380 31260 39432
rect 34612 39380 34664 39432
rect 35808 39380 35860 39432
rect 35992 39491 36044 39500
rect 35992 39457 36001 39491
rect 36001 39457 36035 39491
rect 36035 39457 36044 39491
rect 35992 39448 36044 39457
rect 36912 39380 36964 39432
rect 38292 39448 38344 39500
rect 40408 39448 40460 39500
rect 41144 39448 41196 39500
rect 37372 39380 37424 39432
rect 40224 39380 40276 39432
rect 40684 39380 40736 39432
rect 41604 39423 41656 39432
rect 41604 39389 41613 39423
rect 41613 39389 41647 39423
rect 41647 39389 41656 39423
rect 41604 39380 41656 39389
rect 43076 39491 43128 39500
rect 43076 39457 43085 39491
rect 43085 39457 43119 39491
rect 43119 39457 43128 39491
rect 43076 39448 43128 39457
rect 45376 39584 45428 39636
rect 46204 39516 46256 39568
rect 46664 39627 46716 39636
rect 46664 39593 46673 39627
rect 46673 39593 46707 39627
rect 46707 39593 46716 39627
rect 46664 39584 46716 39593
rect 47400 39627 47452 39636
rect 47400 39593 47409 39627
rect 47409 39593 47443 39627
rect 47443 39593 47452 39627
rect 47400 39584 47452 39593
rect 48412 39627 48464 39636
rect 48412 39593 48421 39627
rect 48421 39593 48455 39627
rect 48455 39593 48464 39627
rect 48412 39584 48464 39593
rect 48596 39584 48648 39636
rect 49608 39516 49660 39568
rect 50528 39627 50580 39636
rect 50528 39593 50537 39627
rect 50537 39593 50571 39627
rect 50571 39593 50580 39627
rect 50528 39584 50580 39593
rect 54576 39584 54628 39636
rect 54944 39584 54996 39636
rect 55312 39627 55364 39636
rect 55312 39593 55321 39627
rect 55321 39593 55355 39627
rect 55355 39593 55364 39627
rect 55312 39584 55364 39593
rect 55956 39584 56008 39636
rect 53748 39559 53800 39568
rect 53748 39525 53757 39559
rect 53757 39525 53791 39559
rect 53791 39525 53800 39559
rect 53748 39516 53800 39525
rect 56508 39516 56560 39568
rect 57244 39516 57296 39568
rect 58440 39584 58492 39636
rect 43444 39380 43496 39432
rect 43812 39380 43864 39432
rect 44548 39380 44600 39432
rect 47492 39423 47544 39432
rect 47492 39389 47501 39423
rect 47501 39389 47535 39423
rect 47535 39389 47544 39423
rect 47492 39380 47544 39389
rect 47768 39380 47820 39432
rect 50620 39491 50672 39500
rect 50620 39457 50629 39491
rect 50629 39457 50663 39491
rect 50663 39457 50672 39491
rect 50620 39448 50672 39457
rect 50804 39448 50856 39500
rect 49516 39380 49568 39432
rect 29368 39244 29420 39296
rect 29460 39244 29512 39296
rect 31392 39244 31444 39296
rect 32680 39244 32732 39296
rect 32772 39244 32824 39296
rect 34336 39244 34388 39296
rect 35072 39244 35124 39296
rect 35440 39287 35492 39296
rect 35440 39253 35449 39287
rect 35449 39253 35483 39287
rect 35483 39253 35492 39287
rect 35440 39244 35492 39253
rect 37372 39244 37424 39296
rect 40132 39244 40184 39296
rect 40592 39244 40644 39296
rect 41052 39287 41104 39296
rect 41052 39253 41061 39287
rect 41061 39253 41095 39287
rect 41095 39253 41104 39287
rect 41052 39244 41104 39253
rect 41788 39244 41840 39296
rect 42432 39244 42484 39296
rect 42616 39287 42668 39296
rect 42616 39253 42625 39287
rect 42625 39253 42659 39287
rect 42659 39253 42668 39287
rect 42616 39244 42668 39253
rect 44824 39287 44876 39296
rect 44824 39253 44833 39287
rect 44833 39253 44867 39287
rect 44867 39253 44876 39287
rect 44824 39244 44876 39253
rect 50160 39423 50212 39432
rect 50160 39389 50169 39423
rect 50169 39389 50203 39423
rect 50203 39389 50212 39423
rect 50160 39380 50212 39389
rect 50528 39380 50580 39432
rect 52552 39448 52604 39500
rect 53656 39448 53708 39500
rect 54484 39423 54536 39432
rect 54484 39389 54493 39423
rect 54493 39389 54527 39423
rect 54527 39389 54536 39423
rect 54484 39380 54536 39389
rect 54576 39423 54628 39432
rect 54576 39389 54585 39423
rect 54585 39389 54619 39423
rect 54619 39389 54628 39423
rect 54576 39380 54628 39389
rect 54852 39380 54904 39432
rect 55036 39380 55088 39432
rect 52736 39244 52788 39296
rect 54208 39312 54260 39364
rect 57152 39423 57204 39432
rect 57152 39389 57161 39423
rect 57161 39389 57195 39423
rect 57195 39389 57204 39423
rect 57152 39380 57204 39389
rect 57336 39423 57388 39432
rect 57336 39389 57345 39423
rect 57345 39389 57379 39423
rect 57379 39389 57388 39423
rect 57336 39380 57388 39389
rect 57704 39380 57756 39432
rect 59268 39380 59320 39432
rect 55220 39244 55272 39296
rect 56140 39244 56192 39296
rect 58808 39312 58860 39364
rect 57796 39244 57848 39296
rect 1998 39142 2050 39194
rect 2062 39142 2114 39194
rect 2126 39142 2178 39194
rect 2190 39142 2242 39194
rect 2254 39142 2306 39194
rect 50998 39142 51050 39194
rect 51062 39142 51114 39194
rect 51126 39142 51178 39194
rect 51190 39142 51242 39194
rect 51254 39142 51306 39194
rect 8208 39083 8260 39092
rect 8208 39049 8217 39083
rect 8217 39049 8251 39083
rect 8251 39049 8260 39083
rect 8208 39040 8260 39049
rect 12532 39040 12584 39092
rect 12256 38972 12308 39024
rect 13820 39040 13872 39092
rect 13912 39040 13964 39092
rect 7104 38904 7156 38956
rect 7932 38904 7984 38956
rect 8392 38904 8444 38956
rect 9312 38904 9364 38956
rect 10324 38947 10376 38956
rect 10324 38913 10333 38947
rect 10333 38913 10367 38947
rect 10367 38913 10376 38947
rect 10324 38904 10376 38913
rect 14004 38972 14056 39024
rect 13176 38947 13228 38956
rect 13176 38913 13185 38947
rect 13185 38913 13219 38947
rect 13219 38913 13228 38947
rect 13176 38904 13228 38913
rect 15108 38904 15160 38956
rect 15384 38947 15436 38956
rect 15384 38913 15393 38947
rect 15393 38913 15427 38947
rect 15427 38913 15436 38947
rect 15384 38904 15436 38913
rect 17500 39040 17552 39092
rect 19340 39040 19392 39092
rect 19708 39040 19760 39092
rect 28954 39040 29006 39092
rect 29276 39083 29328 39092
rect 29276 39049 29306 39083
rect 29306 39049 29328 39083
rect 29276 39040 29328 39049
rect 29644 39040 29696 39092
rect 41788 39040 41840 39092
rect 18512 38972 18564 39024
rect 24124 38972 24176 39024
rect 24676 39015 24728 39024
rect 24676 38981 24685 39015
rect 24685 38981 24719 39015
rect 24719 38981 24728 39015
rect 24676 38972 24728 38981
rect 24952 38972 25004 39024
rect 19892 38947 19944 38956
rect 19892 38913 19901 38947
rect 19901 38913 19935 38947
rect 19935 38913 19944 38947
rect 19892 38904 19944 38913
rect 19984 38947 20036 38956
rect 19984 38913 19993 38947
rect 19993 38913 20027 38947
rect 20027 38913 20036 38947
rect 19984 38904 20036 38913
rect 20628 38904 20680 38956
rect 9680 38836 9732 38888
rect 9956 38836 10008 38888
rect 15568 38836 15620 38888
rect 19432 38836 19484 38888
rect 19616 38836 19668 38888
rect 21364 38904 21416 38956
rect 24492 38947 24544 38956
rect 24492 38913 24501 38947
rect 24501 38913 24535 38947
rect 24535 38913 24544 38947
rect 24492 38904 24544 38913
rect 25136 38947 25188 38956
rect 25136 38913 25145 38947
rect 25145 38913 25179 38947
rect 25179 38913 25188 38947
rect 25136 38904 25188 38913
rect 26240 38904 26292 38956
rect 26884 39015 26936 39024
rect 26884 38981 26893 39015
rect 26893 38981 26927 39015
rect 26927 38981 26936 39015
rect 26884 38972 26936 38981
rect 30840 38972 30892 39024
rect 32220 38972 32272 39024
rect 28908 38904 28960 38956
rect 30012 38904 30064 38956
rect 30564 38904 30616 38956
rect 31116 38904 31168 38956
rect 32128 38904 32180 38956
rect 33692 38972 33744 39024
rect 34060 38972 34112 39024
rect 34612 38972 34664 39024
rect 21088 38836 21140 38888
rect 23480 38836 23532 38888
rect 25044 38879 25096 38888
rect 25044 38845 25053 38879
rect 25053 38845 25087 38879
rect 25087 38845 25096 38879
rect 25044 38836 25096 38845
rect 6920 38700 6972 38752
rect 7012 38700 7064 38752
rect 9864 38700 9916 38752
rect 10232 38768 10284 38820
rect 10324 38768 10376 38820
rect 12072 38811 12124 38820
rect 12072 38777 12081 38811
rect 12081 38777 12115 38811
rect 12115 38777 12124 38811
rect 12072 38768 12124 38777
rect 16212 38768 16264 38820
rect 20536 38768 20588 38820
rect 23204 38768 23256 38820
rect 10968 38700 11020 38752
rect 13820 38700 13872 38752
rect 15384 38700 15436 38752
rect 16396 38700 16448 38752
rect 20260 38743 20312 38752
rect 20260 38709 20269 38743
rect 20269 38709 20303 38743
rect 20303 38709 20312 38743
rect 20260 38700 20312 38709
rect 20352 38700 20404 38752
rect 20720 38700 20772 38752
rect 20812 38700 20864 38752
rect 21824 38700 21876 38752
rect 23020 38743 23072 38752
rect 23020 38709 23029 38743
rect 23029 38709 23063 38743
rect 23063 38709 23072 38743
rect 23020 38700 23072 38709
rect 23756 38700 23808 38752
rect 26148 38879 26200 38888
rect 26148 38845 26157 38879
rect 26157 38845 26191 38879
rect 26191 38845 26200 38879
rect 26148 38836 26200 38845
rect 27620 38836 27672 38888
rect 28540 38836 28592 38888
rect 27804 38768 27856 38820
rect 28632 38768 28684 38820
rect 25688 38700 25740 38752
rect 28954 38700 29006 38752
rect 29092 38700 29144 38752
rect 31576 38768 31628 38820
rect 32772 38811 32824 38820
rect 32772 38777 32781 38811
rect 32781 38777 32815 38811
rect 32815 38777 32824 38811
rect 32772 38768 32824 38777
rect 30840 38743 30892 38752
rect 30840 38709 30849 38743
rect 30849 38709 30883 38743
rect 30883 38709 30892 38743
rect 30840 38700 30892 38709
rect 31208 38743 31260 38752
rect 31208 38709 31217 38743
rect 31217 38709 31251 38743
rect 31251 38709 31260 38743
rect 31208 38700 31260 38709
rect 31392 38700 31444 38752
rect 32128 38700 32180 38752
rect 33968 38904 34020 38956
rect 37188 38904 37240 38956
rect 39120 38972 39172 39024
rect 39304 39015 39356 39024
rect 39304 38981 39313 39015
rect 39313 38981 39347 39015
rect 39347 38981 39356 39015
rect 39304 38972 39356 38981
rect 40132 38972 40184 39024
rect 37372 38947 37424 38956
rect 37372 38913 37381 38947
rect 37381 38913 37415 38947
rect 37415 38913 37424 38947
rect 37372 38904 37424 38913
rect 38200 38904 38252 38956
rect 38292 38947 38344 38956
rect 38292 38913 38301 38947
rect 38301 38913 38335 38947
rect 38335 38913 38344 38947
rect 38292 38904 38344 38913
rect 38476 38904 38528 38956
rect 40224 38904 40276 38956
rect 40592 38947 40644 38956
rect 40592 38913 40601 38947
rect 40601 38913 40635 38947
rect 40635 38913 40644 38947
rect 40592 38904 40644 38913
rect 41236 38904 41288 38956
rect 42892 38904 42944 38956
rect 43444 39040 43496 39092
rect 47492 39040 47544 39092
rect 47676 39083 47728 39092
rect 47676 39049 47685 39083
rect 47685 39049 47719 39083
rect 47719 39049 47728 39083
rect 47676 39040 47728 39049
rect 48320 39040 48372 39092
rect 48964 39040 49016 39092
rect 54208 39083 54260 39092
rect 54208 39049 54217 39083
rect 54217 39049 54251 39083
rect 54251 39049 54260 39083
rect 54208 39040 54260 39049
rect 54484 39040 54536 39092
rect 43628 38972 43680 39024
rect 43996 38904 44048 38956
rect 45560 38904 45612 38956
rect 33968 38768 34020 38820
rect 34152 38768 34204 38820
rect 35624 38811 35676 38820
rect 35624 38777 35633 38811
rect 35633 38777 35667 38811
rect 35667 38777 35676 38811
rect 35624 38768 35676 38777
rect 34336 38700 34388 38752
rect 38936 38836 38988 38888
rect 41052 38836 41104 38888
rect 41880 38836 41932 38888
rect 43352 38836 43404 38888
rect 45284 38836 45336 38888
rect 48320 38947 48372 38956
rect 48320 38913 48329 38947
rect 48329 38913 48363 38947
rect 48363 38913 48372 38947
rect 48320 38904 48372 38913
rect 50344 38972 50396 39024
rect 50620 38972 50672 39024
rect 49332 38947 49384 38956
rect 49332 38913 49341 38947
rect 49341 38913 49375 38947
rect 49375 38913 49384 38947
rect 49332 38904 49384 38913
rect 49792 38904 49844 38956
rect 50804 38904 50856 38956
rect 54576 38972 54628 39024
rect 48412 38836 48464 38888
rect 49516 38836 49568 38888
rect 37004 38700 37056 38752
rect 37464 38700 37516 38752
rect 38016 38700 38068 38752
rect 38200 38700 38252 38752
rect 41696 38768 41748 38820
rect 45192 38768 45244 38820
rect 45468 38811 45520 38820
rect 45468 38777 45477 38811
rect 45477 38777 45511 38811
rect 45511 38777 45520 38811
rect 45468 38768 45520 38777
rect 46204 38811 46256 38820
rect 46204 38777 46213 38811
rect 46213 38777 46247 38811
rect 46247 38777 46256 38811
rect 46204 38768 46256 38777
rect 46664 38768 46716 38820
rect 47492 38768 47544 38820
rect 49700 38768 49752 38820
rect 50528 38836 50580 38888
rect 52460 38947 52512 38956
rect 52460 38913 52469 38947
rect 52469 38913 52503 38947
rect 52503 38913 52512 38947
rect 52460 38904 52512 38913
rect 53472 38904 53524 38956
rect 55220 38947 55272 38956
rect 55220 38913 55229 38947
rect 55229 38913 55263 38947
rect 55263 38913 55272 38947
rect 55220 38904 55272 38913
rect 55680 38904 55732 38956
rect 58072 39040 58124 39092
rect 58808 39083 58860 39092
rect 58808 39049 58817 39083
rect 58817 39049 58851 39083
rect 58851 39049 58860 39083
rect 58808 39040 58860 39049
rect 58900 39083 58952 39092
rect 58900 39049 58909 39083
rect 58909 39049 58943 39083
rect 58943 39049 58952 39083
rect 58900 39040 58952 39049
rect 52276 38879 52328 38888
rect 52276 38845 52285 38879
rect 52285 38845 52319 38879
rect 52319 38845 52328 38879
rect 52276 38836 52328 38845
rect 53840 38836 53892 38888
rect 55128 38836 55180 38888
rect 55956 38836 56008 38888
rect 50712 38768 50764 38820
rect 52736 38811 52788 38820
rect 52736 38777 52745 38811
rect 52745 38777 52779 38811
rect 52779 38777 52788 38811
rect 52736 38768 52788 38777
rect 56508 38904 56560 38956
rect 57980 38904 58032 38956
rect 59452 38947 59504 38956
rect 59452 38913 59461 38947
rect 59461 38913 59495 38947
rect 59495 38913 59504 38947
rect 59452 38904 59504 38913
rect 56140 38879 56192 38888
rect 56140 38845 56149 38879
rect 56149 38845 56183 38879
rect 56183 38845 56192 38879
rect 56140 38836 56192 38845
rect 59268 38879 59320 38888
rect 59268 38845 59277 38879
rect 59277 38845 59311 38879
rect 59311 38845 59320 38879
rect 59268 38836 59320 38845
rect 39672 38743 39724 38752
rect 39672 38709 39681 38743
rect 39681 38709 39715 38743
rect 39715 38709 39724 38743
rect 39672 38700 39724 38709
rect 39856 38700 39908 38752
rect 41512 38743 41564 38752
rect 41512 38709 41521 38743
rect 41521 38709 41555 38743
rect 41555 38709 41564 38743
rect 41512 38700 41564 38709
rect 42248 38700 42300 38752
rect 44180 38700 44232 38752
rect 45376 38743 45428 38752
rect 45376 38709 45385 38743
rect 45385 38709 45419 38743
rect 45419 38709 45428 38743
rect 45376 38700 45428 38709
rect 45560 38700 45612 38752
rect 47124 38700 47176 38752
rect 47768 38743 47820 38752
rect 47768 38709 47777 38743
rect 47777 38709 47811 38743
rect 47811 38709 47820 38743
rect 47768 38700 47820 38709
rect 48964 38700 49016 38752
rect 50988 38700 51040 38752
rect 54116 38700 54168 38752
rect 55128 38743 55180 38752
rect 55128 38709 55137 38743
rect 55137 38709 55171 38743
rect 55171 38709 55180 38743
rect 55128 38700 55180 38709
rect 55772 38743 55824 38752
rect 55772 38709 55781 38743
rect 55781 38709 55815 38743
rect 55815 38709 55824 38743
rect 55772 38700 55824 38709
rect 56232 38743 56284 38752
rect 56232 38709 56241 38743
rect 56241 38709 56275 38743
rect 56275 38709 56284 38743
rect 56232 38700 56284 38709
rect 58348 38768 58400 38820
rect 63684 38768 63736 38820
rect 59268 38700 59320 38752
rect 2918 38598 2970 38650
rect 2982 38598 3034 38650
rect 3046 38598 3098 38650
rect 3110 38598 3162 38650
rect 3174 38598 3226 38650
rect 51918 38598 51970 38650
rect 51982 38598 52034 38650
rect 52046 38598 52098 38650
rect 52110 38598 52162 38650
rect 52174 38598 52226 38650
rect 6920 38539 6972 38548
rect 6920 38505 6929 38539
rect 6929 38505 6963 38539
rect 6963 38505 6972 38539
rect 6920 38496 6972 38505
rect 7840 38496 7892 38548
rect 8208 38496 8260 38548
rect 7380 38335 7432 38344
rect 7380 38301 7389 38335
rect 7389 38301 7423 38335
rect 7423 38301 7432 38335
rect 7380 38292 7432 38301
rect 8392 38360 8444 38412
rect 8484 38360 8536 38412
rect 8760 38496 8812 38548
rect 10968 38539 11020 38548
rect 10968 38505 10977 38539
rect 10977 38505 11011 38539
rect 11011 38505 11020 38539
rect 10968 38496 11020 38505
rect 11060 38496 11112 38548
rect 10232 38428 10284 38480
rect 15200 38496 15252 38548
rect 15568 38496 15620 38548
rect 9956 38360 10008 38412
rect 10324 38360 10376 38412
rect 7932 38335 7984 38344
rect 7932 38301 7941 38335
rect 7941 38301 7975 38335
rect 7975 38301 7984 38335
rect 7932 38292 7984 38301
rect 9956 38224 10008 38276
rect 11428 38360 11480 38412
rect 12072 38403 12124 38412
rect 12072 38369 12081 38403
rect 12081 38369 12115 38403
rect 12115 38369 12124 38403
rect 12072 38360 12124 38369
rect 12716 38360 12768 38412
rect 14280 38428 14332 38480
rect 11520 38335 11572 38344
rect 11520 38301 11529 38335
rect 11529 38301 11563 38335
rect 11563 38301 11572 38335
rect 11520 38292 11572 38301
rect 12164 38335 12216 38344
rect 12164 38301 12173 38335
rect 12173 38301 12207 38335
rect 12207 38301 12216 38335
rect 12164 38292 12216 38301
rect 12256 38335 12308 38344
rect 12256 38301 12265 38335
rect 12265 38301 12299 38335
rect 12299 38301 12308 38335
rect 12256 38292 12308 38301
rect 11612 38224 11664 38276
rect 12440 38224 12492 38276
rect 12808 38335 12860 38344
rect 12808 38301 12817 38335
rect 12817 38301 12851 38335
rect 12851 38301 12860 38335
rect 12808 38292 12860 38301
rect 15292 38292 15344 38344
rect 16212 38428 16264 38480
rect 14648 38224 14700 38276
rect 14004 38156 14056 38208
rect 15108 38199 15160 38208
rect 15108 38165 15117 38199
rect 15117 38165 15151 38199
rect 15151 38165 15160 38199
rect 15108 38156 15160 38165
rect 16396 38292 16448 38344
rect 17224 38403 17276 38412
rect 17224 38369 17233 38403
rect 17233 38369 17267 38403
rect 17267 38369 17276 38403
rect 17224 38360 17276 38369
rect 18144 38428 18196 38480
rect 20444 38496 20496 38548
rect 20904 38496 20956 38548
rect 21088 38539 21140 38548
rect 21088 38505 21097 38539
rect 21097 38505 21131 38539
rect 21131 38505 21140 38539
rect 21088 38496 21140 38505
rect 23480 38496 23532 38548
rect 23756 38428 23808 38480
rect 21548 38403 21600 38412
rect 21548 38369 21557 38403
rect 21557 38369 21591 38403
rect 21591 38369 21600 38403
rect 21548 38360 21600 38369
rect 25136 38539 25188 38548
rect 25136 38505 25145 38539
rect 25145 38505 25179 38539
rect 25179 38505 25188 38539
rect 25136 38496 25188 38505
rect 26056 38496 26108 38548
rect 27528 38496 27580 38548
rect 27620 38496 27672 38548
rect 34428 38496 34480 38548
rect 34520 38496 34572 38548
rect 29828 38428 29880 38480
rect 25412 38360 25464 38412
rect 30564 38428 30616 38480
rect 30748 38428 30800 38480
rect 33968 38428 34020 38480
rect 35440 38539 35492 38548
rect 35440 38505 35449 38539
rect 35449 38505 35483 38539
rect 35483 38505 35492 38539
rect 35440 38496 35492 38505
rect 35624 38496 35676 38548
rect 38476 38539 38528 38548
rect 38476 38505 38485 38539
rect 38485 38505 38519 38539
rect 38519 38505 38528 38539
rect 38476 38496 38528 38505
rect 37004 38471 37056 38480
rect 37004 38437 37013 38471
rect 37013 38437 37047 38471
rect 37047 38437 37056 38471
rect 37004 38428 37056 38437
rect 30472 38403 30524 38412
rect 30472 38369 30481 38403
rect 30481 38369 30515 38403
rect 30515 38369 30524 38403
rect 30472 38360 30524 38369
rect 17684 38335 17736 38344
rect 17684 38301 17693 38335
rect 17693 38301 17727 38335
rect 17727 38301 17736 38335
rect 17684 38292 17736 38301
rect 19340 38335 19392 38344
rect 19340 38301 19349 38335
rect 19349 38301 19383 38335
rect 19383 38301 19392 38335
rect 19340 38292 19392 38301
rect 20260 38292 20312 38344
rect 22836 38292 22888 38344
rect 23664 38292 23716 38344
rect 26148 38292 26200 38344
rect 26884 38335 26936 38344
rect 26884 38301 26893 38335
rect 26893 38301 26927 38335
rect 26927 38301 26936 38335
rect 26884 38292 26936 38301
rect 16120 38199 16172 38208
rect 16120 38165 16129 38199
rect 16129 38165 16163 38199
rect 16163 38165 16172 38199
rect 16120 38156 16172 38165
rect 26240 38224 26292 38276
rect 19064 38156 19116 38208
rect 19248 38156 19300 38208
rect 23480 38156 23532 38208
rect 25688 38156 25740 38208
rect 26792 38224 26844 38276
rect 27804 38335 27856 38344
rect 27804 38301 27813 38335
rect 27813 38301 27847 38335
rect 27847 38301 27856 38335
rect 27804 38292 27856 38301
rect 29184 38292 29236 38344
rect 28172 38224 28224 38276
rect 28632 38156 28684 38208
rect 30012 38292 30064 38344
rect 31392 38360 31444 38412
rect 33140 38360 33192 38412
rect 31116 38335 31168 38344
rect 31116 38301 31125 38335
rect 31125 38301 31159 38335
rect 31159 38301 31168 38335
rect 31116 38292 31168 38301
rect 31484 38292 31536 38344
rect 34244 38292 34296 38344
rect 34704 38292 34756 38344
rect 36728 38403 36780 38412
rect 36728 38369 36737 38403
rect 36737 38369 36771 38403
rect 36771 38369 36780 38403
rect 36728 38360 36780 38369
rect 40868 38496 40920 38548
rect 41420 38496 41472 38548
rect 42616 38496 42668 38548
rect 42708 38496 42760 38548
rect 39856 38428 39908 38480
rect 40040 38428 40092 38480
rect 44548 38428 44600 38480
rect 45192 38496 45244 38548
rect 46204 38496 46256 38548
rect 47768 38496 47820 38548
rect 48964 38471 49016 38480
rect 48964 38437 48973 38471
rect 48973 38437 49007 38471
rect 49007 38437 49016 38471
rect 48964 38428 49016 38437
rect 49700 38428 49752 38480
rect 50344 38496 50396 38548
rect 50988 38539 51040 38548
rect 50988 38505 50997 38539
rect 50997 38505 51031 38539
rect 51031 38505 51040 38539
rect 50988 38496 51040 38505
rect 63776 38496 63828 38548
rect 53840 38428 53892 38480
rect 55772 38428 55824 38480
rect 55956 38428 56008 38480
rect 58348 38428 58400 38480
rect 60740 38428 60792 38480
rect 62488 38428 62540 38480
rect 35164 38335 35216 38344
rect 35164 38301 35173 38335
rect 35173 38301 35207 38335
rect 35207 38301 35216 38335
rect 35164 38292 35216 38301
rect 35256 38292 35308 38344
rect 40868 38360 40920 38412
rect 41328 38360 41380 38412
rect 43260 38403 43312 38412
rect 43260 38369 43269 38403
rect 43269 38369 43303 38403
rect 43303 38369 43312 38403
rect 43260 38360 43312 38369
rect 45284 38403 45336 38412
rect 45284 38369 45293 38403
rect 45293 38369 45327 38403
rect 45327 38369 45336 38403
rect 45284 38360 45336 38369
rect 38752 38292 38804 38344
rect 39948 38292 40000 38344
rect 40776 38292 40828 38344
rect 41604 38292 41656 38344
rect 42524 38335 42576 38344
rect 42524 38301 42533 38335
rect 42533 38301 42567 38335
rect 42567 38301 42576 38335
rect 42524 38292 42576 38301
rect 44456 38292 44508 38344
rect 29552 38224 29604 38276
rect 30656 38199 30708 38208
rect 30656 38165 30665 38199
rect 30665 38165 30699 38199
rect 30699 38165 30708 38199
rect 30656 38156 30708 38165
rect 32220 38199 32272 38208
rect 32220 38165 32229 38199
rect 32229 38165 32263 38199
rect 32263 38165 32272 38199
rect 32220 38156 32272 38165
rect 41512 38224 41564 38276
rect 40776 38156 40828 38208
rect 41328 38156 41380 38208
rect 43996 38224 44048 38276
rect 43812 38156 43864 38208
rect 44824 38156 44876 38208
rect 46572 38335 46624 38344
rect 46572 38301 46581 38335
rect 46581 38301 46615 38335
rect 46615 38301 46624 38335
rect 46572 38292 46624 38301
rect 47308 38360 47360 38412
rect 47676 38360 47728 38412
rect 48228 38360 48280 38412
rect 50804 38360 50856 38412
rect 46756 38292 46808 38344
rect 50896 38292 50948 38344
rect 51724 38292 51776 38344
rect 49976 38224 50028 38276
rect 54116 38292 54168 38344
rect 54392 38292 54444 38344
rect 55220 38335 55272 38344
rect 55220 38301 55229 38335
rect 55229 38301 55263 38335
rect 55263 38301 55272 38335
rect 55220 38292 55272 38301
rect 57796 38335 57848 38344
rect 57796 38301 57805 38335
rect 57805 38301 57839 38335
rect 57839 38301 57848 38335
rect 57796 38292 57848 38301
rect 58164 38292 58216 38344
rect 58440 38292 58492 38344
rect 64972 38360 65024 38412
rect 59268 38292 59320 38344
rect 56784 38224 56836 38276
rect 47492 38156 47544 38208
rect 50620 38199 50672 38208
rect 50620 38165 50629 38199
rect 50629 38165 50663 38199
rect 50663 38165 50672 38199
rect 50620 38156 50672 38165
rect 51632 38156 51684 38208
rect 57152 38156 57204 38208
rect 57704 38156 57756 38208
rect 63316 38156 63368 38208
rect 1998 38054 2050 38106
rect 2062 38054 2114 38106
rect 2126 38054 2178 38106
rect 2190 38054 2242 38106
rect 2254 38054 2306 38106
rect 50998 38054 51050 38106
rect 51062 38054 51114 38106
rect 51126 38054 51178 38106
rect 51190 38054 51242 38106
rect 51254 38054 51306 38106
rect 7380 37952 7432 38004
rect 9864 37952 9916 38004
rect 15384 37952 15436 38004
rect 16120 37952 16172 38004
rect 17224 37995 17276 38004
rect 17224 37961 17233 37995
rect 17233 37961 17267 37995
rect 17267 37961 17276 37995
rect 17224 37952 17276 37961
rect 19340 37952 19392 38004
rect 7932 37884 7984 37936
rect 7104 37816 7156 37868
rect 12440 37884 12492 37936
rect 14648 37884 14700 37936
rect 18052 37884 18104 37936
rect 22836 37884 22888 37936
rect 23296 37884 23348 37936
rect 12256 37816 12308 37868
rect 12808 37816 12860 37868
rect 15108 37816 15160 37868
rect 15200 37816 15252 37868
rect 11520 37748 11572 37800
rect 14280 37748 14332 37800
rect 16212 37791 16264 37800
rect 16212 37757 16221 37791
rect 16221 37757 16255 37791
rect 16255 37757 16264 37791
rect 16212 37748 16264 37757
rect 18696 37748 18748 37800
rect 19156 37791 19208 37800
rect 19156 37757 19165 37791
rect 19165 37757 19199 37791
rect 19199 37757 19208 37791
rect 19156 37748 19208 37757
rect 7012 37680 7064 37732
rect 9036 37680 9088 37732
rect 8760 37655 8812 37664
rect 8760 37621 8769 37655
rect 8769 37621 8803 37655
rect 8803 37621 8812 37655
rect 8760 37612 8812 37621
rect 9956 37655 10008 37664
rect 9956 37621 9965 37655
rect 9965 37621 9999 37655
rect 9999 37621 10008 37655
rect 9956 37612 10008 37621
rect 12072 37680 12124 37732
rect 19248 37680 19300 37732
rect 23388 37816 23440 37868
rect 25688 37952 25740 38004
rect 26884 37952 26936 38004
rect 23020 37748 23072 37800
rect 20720 37680 20772 37732
rect 20812 37723 20864 37732
rect 20812 37689 20821 37723
rect 20821 37689 20855 37723
rect 20855 37689 20864 37723
rect 20812 37680 20864 37689
rect 20904 37680 20956 37732
rect 10508 37612 10560 37664
rect 15016 37612 15068 37664
rect 22284 37655 22336 37664
rect 22284 37621 22293 37655
rect 22293 37621 22327 37655
rect 22327 37621 22336 37655
rect 22284 37612 22336 37621
rect 23848 37612 23900 37664
rect 25412 37680 25464 37732
rect 26148 37816 26200 37868
rect 27620 37884 27672 37936
rect 27988 37884 28040 37936
rect 28632 37859 28684 37868
rect 28632 37825 28641 37859
rect 28641 37825 28675 37859
rect 28675 37825 28684 37859
rect 28632 37816 28684 37825
rect 30656 37884 30708 37936
rect 30288 37816 30340 37868
rect 27620 37748 27672 37800
rect 27896 37748 27948 37800
rect 32036 37859 32088 37868
rect 32036 37825 32045 37859
rect 32045 37825 32079 37859
rect 32079 37825 32088 37859
rect 32036 37816 32088 37825
rect 30656 37748 30708 37800
rect 26516 37723 26568 37732
rect 26516 37689 26525 37723
rect 26525 37689 26559 37723
rect 26559 37689 26568 37723
rect 26516 37680 26568 37689
rect 27804 37612 27856 37664
rect 29184 37680 29236 37732
rect 28540 37655 28592 37664
rect 28540 37621 28549 37655
rect 28549 37621 28583 37655
rect 28583 37621 28592 37655
rect 28540 37612 28592 37621
rect 29644 37612 29696 37664
rect 30012 37612 30064 37664
rect 31668 37680 31720 37732
rect 31852 37680 31904 37732
rect 34244 37927 34296 37936
rect 34244 37893 34253 37927
rect 34253 37893 34287 37927
rect 34287 37893 34296 37927
rect 34244 37884 34296 37893
rect 34336 37884 34388 37936
rect 35164 37816 35216 37868
rect 37096 37859 37148 37868
rect 37096 37825 37105 37859
rect 37105 37825 37139 37859
rect 37139 37825 37148 37859
rect 37096 37816 37148 37825
rect 37188 37859 37240 37868
rect 37188 37825 37197 37859
rect 37197 37825 37231 37859
rect 37231 37825 37240 37859
rect 37188 37816 37240 37825
rect 38936 37927 38988 37936
rect 38936 37893 38945 37927
rect 38945 37893 38979 37927
rect 38979 37893 38988 37927
rect 38936 37884 38988 37893
rect 39948 37884 40000 37936
rect 35348 37791 35400 37800
rect 35348 37757 35357 37791
rect 35357 37757 35391 37791
rect 35391 37757 35400 37791
rect 35348 37748 35400 37757
rect 38752 37748 38804 37800
rect 33784 37612 33836 37664
rect 34336 37612 34388 37664
rect 34520 37612 34572 37664
rect 35440 37612 35492 37664
rect 37464 37723 37516 37732
rect 37464 37689 37473 37723
rect 37473 37689 37507 37723
rect 37507 37689 37516 37723
rect 37464 37680 37516 37689
rect 39948 37612 40000 37664
rect 40408 37859 40460 37868
rect 40408 37825 40417 37859
rect 40417 37825 40451 37859
rect 40451 37825 40460 37859
rect 40408 37816 40460 37825
rect 41052 37816 41104 37868
rect 41144 37816 41196 37868
rect 41328 37816 41380 37868
rect 42708 37884 42760 37936
rect 44180 37995 44232 38004
rect 44180 37961 44189 37995
rect 44189 37961 44223 37995
rect 44223 37961 44232 37995
rect 44180 37952 44232 37961
rect 44456 37995 44508 38004
rect 44456 37961 44465 37995
rect 44465 37961 44499 37995
rect 44499 37961 44508 37995
rect 44456 37952 44508 37961
rect 46756 37952 46808 38004
rect 49976 37952 50028 38004
rect 50620 37952 50672 38004
rect 50712 37952 50764 38004
rect 51724 37995 51776 38004
rect 51724 37961 51733 37995
rect 51733 37961 51767 37995
rect 51767 37961 51776 37995
rect 51724 37952 51776 37961
rect 54392 37995 54444 38004
rect 54392 37961 54401 37995
rect 54401 37961 54435 37995
rect 54435 37961 54444 37995
rect 54392 37952 54444 37961
rect 56232 37952 56284 38004
rect 57888 37952 57940 38004
rect 63868 37952 63920 38004
rect 44088 37816 44140 37868
rect 45008 37859 45060 37868
rect 45008 37825 45017 37859
rect 45017 37825 45051 37859
rect 45051 37825 45060 37859
rect 45008 37816 45060 37825
rect 47124 37816 47176 37868
rect 47860 37816 47912 37868
rect 49700 37816 49752 37868
rect 42248 37748 42300 37800
rect 44824 37791 44876 37800
rect 44824 37757 44833 37791
rect 44833 37757 44867 37791
rect 44867 37757 44876 37791
rect 44824 37748 44876 37757
rect 50160 37816 50212 37868
rect 53840 37884 53892 37936
rect 40960 37680 41012 37732
rect 41144 37680 41196 37732
rect 44548 37680 44600 37732
rect 47860 37723 47912 37732
rect 47860 37689 47869 37723
rect 47869 37689 47903 37723
rect 47903 37689 47912 37723
rect 47860 37680 47912 37689
rect 48320 37680 48372 37732
rect 54852 37816 54904 37868
rect 56600 37884 56652 37936
rect 58440 37884 58492 37936
rect 53472 37791 53524 37800
rect 53472 37757 53481 37791
rect 53481 37757 53515 37791
rect 53515 37757 53524 37791
rect 53472 37748 53524 37757
rect 55220 37748 55272 37800
rect 53196 37723 53248 37732
rect 53196 37689 53205 37723
rect 53205 37689 53239 37723
rect 53239 37689 53248 37723
rect 53196 37680 53248 37689
rect 53932 37723 53984 37732
rect 53932 37689 53941 37723
rect 53941 37689 53975 37723
rect 53975 37689 53984 37723
rect 53932 37680 53984 37689
rect 54208 37680 54260 37732
rect 55128 37680 55180 37732
rect 55404 37723 55456 37732
rect 55404 37689 55413 37723
rect 55413 37689 55447 37723
rect 55447 37689 55456 37723
rect 55404 37680 55456 37689
rect 42064 37612 42116 37664
rect 43812 37655 43864 37664
rect 43812 37621 43821 37655
rect 43821 37621 43855 37655
rect 43855 37621 43864 37655
rect 43812 37612 43864 37621
rect 45376 37612 45428 37664
rect 47584 37612 47636 37664
rect 48412 37612 48464 37664
rect 51724 37612 51776 37664
rect 51816 37612 51868 37664
rect 57888 37859 57940 37868
rect 57888 37825 57897 37859
rect 57897 37825 57931 37859
rect 57931 37825 57940 37859
rect 57888 37816 57940 37825
rect 57980 37816 58032 37868
rect 63132 37816 63184 37868
rect 63684 37859 63736 37868
rect 63684 37825 63693 37859
rect 63693 37825 63727 37859
rect 63727 37825 63736 37859
rect 63684 37816 63736 37825
rect 63776 37859 63828 37868
rect 63776 37825 63785 37859
rect 63785 37825 63819 37859
rect 63819 37825 63828 37859
rect 63776 37816 63828 37825
rect 58348 37748 58400 37800
rect 55864 37723 55916 37732
rect 55864 37689 55873 37723
rect 55873 37689 55907 37723
rect 55907 37689 55916 37723
rect 55864 37680 55916 37689
rect 55956 37680 56008 37732
rect 57336 37680 57388 37732
rect 59820 37680 59872 37732
rect 57796 37612 57848 37664
rect 58532 37612 58584 37664
rect 60004 37748 60056 37800
rect 66444 37748 66496 37800
rect 65984 37680 66036 37732
rect 60280 37612 60332 37664
rect 64236 37655 64288 37664
rect 64236 37621 64245 37655
rect 64245 37621 64279 37655
rect 64279 37621 64288 37655
rect 64236 37612 64288 37621
rect 2918 37510 2970 37562
rect 2982 37510 3034 37562
rect 3046 37510 3098 37562
rect 3110 37510 3162 37562
rect 3174 37510 3226 37562
rect 51918 37510 51970 37562
rect 51982 37510 52034 37562
rect 52046 37510 52098 37562
rect 52110 37510 52162 37562
rect 52174 37510 52226 37562
rect 65258 37510 65310 37562
rect 65322 37510 65374 37562
rect 65386 37510 65438 37562
rect 65450 37510 65502 37562
rect 65514 37510 65566 37562
rect 8760 37383 8812 37392
rect 8760 37349 8769 37383
rect 8769 37349 8803 37383
rect 8803 37349 8812 37383
rect 8760 37340 8812 37349
rect 9036 37340 9088 37392
rect 13544 37408 13596 37460
rect 14280 37340 14332 37392
rect 17224 37408 17276 37460
rect 17684 37408 17736 37460
rect 8484 37315 8536 37324
rect 8484 37281 8493 37315
rect 8493 37281 8527 37315
rect 8527 37281 8536 37315
rect 8484 37272 8536 37281
rect 10508 37315 10560 37324
rect 10508 37281 10517 37315
rect 10517 37281 10551 37315
rect 10551 37281 10560 37315
rect 10508 37272 10560 37281
rect 13544 37315 13596 37324
rect 13544 37281 13553 37315
rect 13553 37281 13587 37315
rect 13587 37281 13596 37315
rect 13544 37272 13596 37281
rect 18144 37340 18196 37392
rect 19432 37408 19484 37460
rect 20628 37408 20680 37460
rect 21824 37451 21876 37460
rect 21824 37417 21833 37451
rect 21833 37417 21867 37451
rect 21867 37417 21876 37451
rect 21824 37408 21876 37417
rect 23848 37451 23900 37460
rect 23848 37417 23857 37451
rect 23857 37417 23891 37451
rect 23891 37417 23900 37451
rect 23848 37408 23900 37417
rect 25136 37408 25188 37460
rect 26516 37408 26568 37460
rect 27804 37408 27856 37460
rect 29184 37408 29236 37460
rect 29920 37408 29972 37460
rect 19248 37340 19300 37392
rect 29000 37340 29052 37392
rect 13820 37247 13872 37256
rect 13820 37213 13829 37247
rect 13829 37213 13863 37247
rect 13863 37213 13872 37247
rect 13820 37204 13872 37213
rect 15292 37247 15344 37256
rect 15292 37213 15301 37247
rect 15301 37213 15335 37247
rect 15335 37213 15344 37247
rect 15292 37204 15344 37213
rect 16856 37247 16908 37256
rect 16856 37213 16865 37247
rect 16865 37213 16899 37247
rect 16899 37213 16908 37247
rect 16856 37204 16908 37213
rect 21824 37272 21876 37324
rect 22284 37272 22336 37324
rect 24308 37315 24360 37324
rect 24308 37281 24317 37315
rect 24317 37281 24351 37315
rect 24351 37281 24360 37315
rect 24308 37272 24360 37281
rect 29644 37383 29696 37392
rect 29644 37349 29653 37383
rect 29653 37349 29687 37383
rect 29687 37349 29696 37383
rect 29644 37340 29696 37349
rect 30656 37340 30708 37392
rect 29368 37315 29420 37324
rect 29368 37281 29377 37315
rect 29377 37281 29411 37315
rect 29411 37281 29420 37315
rect 29368 37272 29420 37281
rect 31668 37408 31720 37460
rect 31852 37408 31904 37460
rect 32220 37408 32272 37460
rect 32588 37408 32640 37460
rect 34428 37408 34480 37460
rect 34520 37451 34572 37460
rect 34520 37417 34529 37451
rect 34529 37417 34563 37451
rect 34563 37417 34572 37451
rect 34520 37408 34572 37417
rect 35256 37408 35308 37460
rect 35440 37451 35492 37460
rect 35440 37417 35449 37451
rect 35449 37417 35483 37451
rect 35483 37417 35492 37451
rect 35440 37408 35492 37417
rect 35808 37451 35860 37460
rect 35808 37417 35817 37451
rect 35817 37417 35851 37451
rect 35851 37417 35860 37451
rect 35808 37408 35860 37417
rect 36636 37408 36688 37460
rect 38752 37408 38804 37460
rect 39120 37408 39172 37460
rect 40776 37408 40828 37460
rect 31760 37340 31812 37392
rect 31852 37272 31904 37324
rect 31944 37272 31996 37324
rect 18880 37204 18932 37256
rect 20720 37204 20772 37256
rect 21916 37204 21968 37256
rect 26240 37204 26292 37256
rect 27436 37247 27488 37256
rect 27436 37213 27445 37247
rect 27445 37213 27479 37247
rect 27479 37213 27488 37247
rect 27436 37204 27488 37213
rect 32036 37204 32088 37256
rect 27620 37068 27672 37120
rect 33784 37136 33836 37188
rect 31484 37068 31536 37120
rect 34520 37272 34572 37324
rect 40960 37451 41012 37460
rect 40960 37417 40969 37451
rect 40969 37417 41003 37451
rect 41003 37417 41012 37451
rect 40960 37408 41012 37417
rect 46572 37408 46624 37460
rect 47492 37451 47544 37460
rect 47492 37417 47501 37451
rect 47501 37417 47535 37451
rect 47535 37417 47544 37451
rect 47492 37408 47544 37417
rect 47860 37451 47912 37460
rect 47860 37417 47869 37451
rect 47869 37417 47903 37451
rect 47903 37417 47912 37451
rect 47860 37408 47912 37417
rect 50068 37408 50120 37460
rect 50712 37408 50764 37460
rect 50896 37408 50948 37460
rect 34704 37204 34756 37256
rect 36912 37272 36964 37324
rect 36084 37247 36136 37256
rect 36084 37213 36093 37247
rect 36093 37213 36127 37247
rect 36127 37213 36136 37247
rect 36084 37204 36136 37213
rect 38568 37204 38620 37256
rect 38936 37272 38988 37324
rect 39948 37272 40000 37324
rect 41328 37315 41380 37324
rect 41328 37281 41337 37315
rect 41337 37281 41371 37315
rect 41371 37281 41380 37315
rect 41328 37272 41380 37281
rect 42064 37272 42116 37324
rect 46756 37340 46808 37392
rect 47584 37340 47636 37392
rect 50068 37272 50120 37324
rect 51632 37383 51684 37392
rect 51632 37349 51641 37383
rect 51641 37349 51675 37383
rect 51675 37349 51684 37383
rect 51632 37340 51684 37349
rect 51724 37340 51776 37392
rect 52276 37340 52328 37392
rect 51816 37272 51868 37324
rect 39672 37136 39724 37188
rect 34980 37068 35032 37120
rect 36084 37068 36136 37120
rect 36176 37068 36228 37120
rect 40868 37204 40920 37256
rect 41236 37204 41288 37256
rect 47124 37204 47176 37256
rect 47308 37247 47360 37256
rect 47308 37213 47317 37247
rect 47317 37213 47351 37247
rect 47351 37213 47360 37247
rect 47308 37204 47360 37213
rect 49700 37204 49752 37256
rect 50528 37247 50580 37256
rect 50528 37213 50537 37247
rect 50537 37213 50571 37247
rect 50571 37213 50580 37247
rect 50528 37204 50580 37213
rect 51448 37247 51500 37256
rect 51448 37213 51457 37247
rect 51457 37213 51491 37247
rect 51491 37213 51500 37247
rect 51448 37204 51500 37213
rect 40040 37136 40092 37188
rect 53196 37272 53248 37324
rect 56784 37408 56836 37460
rect 57336 37451 57388 37460
rect 57336 37417 57345 37451
rect 57345 37417 57379 37451
rect 57379 37417 57388 37451
rect 57336 37408 57388 37417
rect 57704 37451 57756 37460
rect 57704 37417 57713 37451
rect 57713 37417 57747 37451
rect 57747 37417 57756 37451
rect 57704 37408 57756 37417
rect 57796 37451 57848 37460
rect 57796 37417 57805 37451
rect 57805 37417 57839 37451
rect 57839 37417 57848 37451
rect 57796 37408 57848 37417
rect 58164 37451 58216 37460
rect 58164 37417 58173 37451
rect 58173 37417 58207 37451
rect 58207 37417 58216 37451
rect 58164 37408 58216 37417
rect 58532 37451 58584 37460
rect 58532 37417 58541 37451
rect 58541 37417 58575 37451
rect 58575 37417 58584 37451
rect 58532 37408 58584 37417
rect 58624 37451 58676 37460
rect 58624 37417 58633 37451
rect 58633 37417 58667 37451
rect 58667 37417 58676 37451
rect 58624 37408 58676 37417
rect 59268 37408 59320 37460
rect 59728 37451 59780 37460
rect 59728 37417 59737 37451
rect 59737 37417 59771 37451
rect 59771 37417 59780 37451
rect 59728 37408 59780 37417
rect 59820 37408 59872 37460
rect 60280 37451 60332 37460
rect 60280 37417 60289 37451
rect 60289 37417 60323 37451
rect 60323 37417 60332 37451
rect 60280 37408 60332 37417
rect 65156 37408 65208 37460
rect 53656 37272 53708 37324
rect 55220 37340 55272 37392
rect 56416 37340 56468 37392
rect 53564 37247 53616 37256
rect 53564 37213 53573 37247
rect 53573 37213 53607 37247
rect 53607 37213 53616 37247
rect 53564 37204 53616 37213
rect 62764 37340 62816 37392
rect 64972 37340 65024 37392
rect 65708 37340 65760 37392
rect 57796 37272 57848 37324
rect 59912 37272 59964 37324
rect 63132 37315 63184 37324
rect 63132 37281 63141 37315
rect 63141 37281 63175 37315
rect 63175 37281 63184 37315
rect 63132 37272 63184 37281
rect 65156 37272 65208 37324
rect 54852 37204 54904 37256
rect 58716 37247 58768 37256
rect 58716 37213 58725 37247
rect 58725 37213 58759 37247
rect 58759 37213 58768 37247
rect 58716 37204 58768 37213
rect 56416 37111 56468 37120
rect 56416 37077 56425 37111
rect 56425 37077 56459 37111
rect 56459 37077 56468 37111
rect 56416 37068 56468 37077
rect 56600 37136 56652 37188
rect 57612 37136 57664 37188
rect 60464 37247 60516 37256
rect 60464 37213 60473 37247
rect 60473 37213 60507 37247
rect 60507 37213 60516 37247
rect 60464 37204 60516 37213
rect 63408 37247 63460 37256
rect 63408 37213 63417 37247
rect 63417 37213 63451 37247
rect 63451 37213 63460 37247
rect 63408 37204 63460 37213
rect 59452 37136 59504 37188
rect 62948 37068 63000 37120
rect 64788 37068 64840 37120
rect 64972 37068 65024 37120
rect 1998 36966 2050 37018
rect 2062 36966 2114 37018
rect 2126 36966 2178 37018
rect 2190 36966 2242 37018
rect 2254 36966 2306 37018
rect 50998 36966 51050 37018
rect 51062 36966 51114 37018
rect 51126 36966 51178 37018
rect 51190 36966 51242 37018
rect 51254 36966 51306 37018
rect 64338 36966 64390 37018
rect 64402 36966 64454 37018
rect 64466 36966 64518 37018
rect 64530 36966 64582 37018
rect 64594 36966 64646 37018
rect 10508 36864 10560 36916
rect 24768 36864 24820 36916
rect 31668 36864 31720 36916
rect 31944 36864 31996 36916
rect 51448 36864 51500 36916
rect 54576 36864 54628 36916
rect 63408 36864 63460 36916
rect 25872 36796 25924 36848
rect 35808 36796 35860 36848
rect 38660 36796 38712 36848
rect 19156 36728 19208 36780
rect 38568 36728 38620 36780
rect 38752 36728 38804 36780
rect 60464 36796 60516 36848
rect 14556 36660 14608 36712
rect 38660 36660 38712 36712
rect 63776 36728 63828 36780
rect 64236 36728 64288 36780
rect 64788 36796 64840 36848
rect 65892 36796 65944 36848
rect 64696 36728 64748 36780
rect 65984 36771 66036 36780
rect 65984 36737 65993 36771
rect 65993 36737 66027 36771
rect 66027 36737 66036 36771
rect 65984 36728 66036 36737
rect 22008 36592 22060 36644
rect 30472 36592 30524 36644
rect 34428 36592 34480 36644
rect 37648 36592 37700 36644
rect 63500 36592 63552 36644
rect 64972 36592 65024 36644
rect 66260 36592 66312 36644
rect 30288 36524 30340 36576
rect 60832 36524 60884 36576
rect 65064 36524 65116 36576
rect 26976 36456 27028 36508
rect 28816 36456 28868 36508
rect 30380 36456 30432 36508
rect 37280 36456 37332 36508
rect 33048 36388 33100 36440
rect 65258 36422 65310 36474
rect 65322 36422 65374 36474
rect 65386 36422 65438 36474
rect 65450 36422 65502 36474
rect 65514 36422 65566 36474
rect 21640 36320 21692 36372
rect 42708 36320 42760 36372
rect 65616 36363 65668 36372
rect 65616 36329 65625 36363
rect 65625 36329 65659 36363
rect 65659 36329 65668 36363
rect 65616 36320 65668 36329
rect 65984 36320 66036 36372
rect 23204 36252 23256 36304
rect 63592 36252 63644 36304
rect 65432 36252 65484 36304
rect 65708 36252 65760 36304
rect 20076 35912 20128 35964
rect 28724 36184 28776 36236
rect 28816 36184 28868 36236
rect 33048 36184 33100 36236
rect 42616 36184 42668 36236
rect 59360 36184 59412 36236
rect 23572 36116 23624 36168
rect 62120 36116 62172 36168
rect 63868 36159 63920 36168
rect 63868 36125 63877 36159
rect 63877 36125 63911 36159
rect 63911 36125 63920 36159
rect 63868 36116 63920 36125
rect 64236 36116 64288 36168
rect 24492 36048 24544 36100
rect 63132 36048 63184 36100
rect 25228 35980 25280 36032
rect 64788 35980 64840 36032
rect 24308 35912 24360 35964
rect 21364 35844 21416 35896
rect 24768 35844 24820 35896
rect 30104 35844 30156 35896
rect 36544 35844 36596 35896
rect 64338 35878 64390 35930
rect 64402 35878 64454 35930
rect 64466 35878 64518 35930
rect 64530 35878 64582 35930
rect 64594 35878 64646 35930
rect 27620 35776 27672 35828
rect 64236 35776 64288 35828
rect 8208 35708 8260 35760
rect 14832 35708 14884 35760
rect 59360 35708 59412 35760
rect 65708 35708 65760 35760
rect 22192 35640 22244 35692
rect 42616 35640 42668 35692
rect 63684 35640 63736 35692
rect 65156 35640 65208 35692
rect 65892 35640 65944 35692
rect 66076 35640 66128 35692
rect 23020 35572 23072 35624
rect 62028 35572 62080 35624
rect 65064 35615 65116 35624
rect 65064 35581 65073 35615
rect 65073 35581 65107 35615
rect 65107 35581 65116 35615
rect 65064 35572 65116 35581
rect 60832 35504 60884 35556
rect 63500 35504 63552 35556
rect 64236 35436 64288 35488
rect 65258 35334 65310 35386
rect 65322 35334 65374 35386
rect 65386 35334 65438 35386
rect 65450 35334 65502 35386
rect 65514 35334 65566 35386
rect 65800 35028 65852 35080
rect 66076 35028 66128 35080
rect 62488 34892 62540 34944
rect 64052 34892 64104 34944
rect 65616 34892 65668 34944
rect 65800 34892 65852 34944
rect 64338 34790 64390 34842
rect 64402 34790 64454 34842
rect 64466 34790 64518 34842
rect 64530 34790 64582 34842
rect 64594 34790 64646 34842
rect 63316 34688 63368 34740
rect 65616 34731 65668 34740
rect 65616 34697 65625 34731
rect 65625 34697 65659 34731
rect 65659 34697 65668 34731
rect 65616 34688 65668 34697
rect 63868 34527 63920 34536
rect 63868 34493 63877 34527
rect 63877 34493 63911 34527
rect 63911 34493 63920 34527
rect 63868 34484 63920 34493
rect 64144 34459 64196 34468
rect 64144 34425 64153 34459
rect 64153 34425 64187 34459
rect 64187 34425 64196 34459
rect 64144 34416 64196 34425
rect 65156 34416 65208 34468
rect 65258 34246 65310 34298
rect 65322 34246 65374 34298
rect 65386 34246 65438 34298
rect 65450 34246 65502 34298
rect 65514 34246 65566 34298
rect 64144 34144 64196 34196
rect 65616 34051 65668 34060
rect 65616 34017 65625 34051
rect 65625 34017 65659 34051
rect 65659 34017 65668 34051
rect 65616 34008 65668 34017
rect 64696 33940 64748 33992
rect 64696 33804 64748 33856
rect 64338 33702 64390 33754
rect 64402 33702 64454 33754
rect 64466 33702 64518 33754
rect 64530 33702 64582 33754
rect 64594 33702 64646 33754
rect 65984 33532 66036 33584
rect 66260 33532 66312 33584
rect 64788 33464 64840 33516
rect 65064 33464 65116 33516
rect 65616 33396 65668 33448
rect 65984 33439 66036 33448
rect 65984 33405 65993 33439
rect 65993 33405 66027 33439
rect 66027 33405 66036 33439
rect 65984 33396 66036 33405
rect 66444 33328 66496 33380
rect 65156 33260 65208 33312
rect 65616 33260 65668 33312
rect 62856 33192 62908 33244
rect 63408 33192 63460 33244
rect 65258 33158 65310 33210
rect 65322 33158 65374 33210
rect 65386 33158 65438 33210
rect 65450 33158 65502 33210
rect 65514 33158 65566 33210
rect 66076 32988 66128 33040
rect 63960 32895 64012 32904
rect 63960 32861 63969 32895
rect 63969 32861 64003 32895
rect 64003 32861 64012 32895
rect 63960 32852 64012 32861
rect 64880 32852 64932 32904
rect 65248 32716 65300 32768
rect 65984 32716 66036 32768
rect 64338 32614 64390 32666
rect 64402 32614 64454 32666
rect 64466 32614 64518 32666
rect 64530 32614 64582 32666
rect 64594 32614 64646 32666
rect 64696 32555 64748 32564
rect 64696 32521 64705 32555
rect 64705 32521 64739 32555
rect 64739 32521 64748 32555
rect 64696 32512 64748 32521
rect 64880 32512 64932 32564
rect 65984 32444 66036 32496
rect 66260 32444 66312 32496
rect 65156 32376 65208 32428
rect 65248 32308 65300 32360
rect 65616 32308 65668 32360
rect 64880 32240 64932 32292
rect 65708 32240 65760 32292
rect 65616 32172 65668 32224
rect 65892 32376 65944 32428
rect 65258 32070 65310 32122
rect 65322 32070 65374 32122
rect 65386 32070 65438 32122
rect 65450 32070 65502 32122
rect 65514 32070 65566 32122
rect 63868 31968 63920 32020
rect 64052 31968 64104 32020
rect 64972 31900 65024 31952
rect 63684 31832 63736 31884
rect 63868 31832 63920 31884
rect 64880 31832 64932 31884
rect 64338 31526 64390 31578
rect 64402 31526 64454 31578
rect 64466 31526 64518 31578
rect 64530 31526 64582 31578
rect 64594 31526 64646 31578
rect 65064 31356 65116 31408
rect 64880 31288 64932 31340
rect 65984 31288 66036 31340
rect 66076 31288 66128 31340
rect 65800 31220 65852 31272
rect 65708 31152 65760 31204
rect 65800 31084 65852 31136
rect 62580 30948 62632 31000
rect 63224 30948 63276 31000
rect 65258 30982 65310 31034
rect 65322 30982 65374 31034
rect 65386 30982 65438 31034
rect 65450 30982 65502 31034
rect 65514 30982 65566 31034
rect 65800 30812 65852 30864
rect 63960 30744 64012 30796
rect 64696 30676 64748 30728
rect 65984 30540 66036 30592
rect 64338 30438 64390 30490
rect 64402 30438 64454 30490
rect 64466 30438 64518 30490
rect 64530 30438 64582 30490
rect 64594 30438 64646 30490
rect 64696 30336 64748 30388
rect 65064 30243 65116 30252
rect 65064 30209 65073 30243
rect 65073 30209 65107 30243
rect 65107 30209 65116 30243
rect 65064 30200 65116 30209
rect 65616 30200 65668 30252
rect 65984 30175 66036 30184
rect 65984 30141 65993 30175
rect 65993 30141 66027 30175
rect 66027 30141 66036 30175
rect 65984 30132 66036 30141
rect 65258 29894 65310 29946
rect 65322 29894 65374 29946
rect 65386 29894 65438 29946
rect 65450 29894 65502 29946
rect 65514 29894 65566 29946
rect 65064 29724 65116 29776
rect 65616 29588 65668 29640
rect 65708 29588 65760 29640
rect 64696 29452 64748 29504
rect 64338 29350 64390 29402
rect 64402 29350 64454 29402
rect 64466 29350 64518 29402
rect 64530 29350 64582 29402
rect 64594 29350 64646 29402
rect 64052 29155 64104 29164
rect 64052 29121 64061 29155
rect 64061 29121 64095 29155
rect 64095 29121 64104 29155
rect 64052 29112 64104 29121
rect 64696 29112 64748 29164
rect 65708 29112 65760 29164
rect 65800 28976 65852 29028
rect 66168 28976 66220 29028
rect 65258 28806 65310 28858
rect 65322 28806 65374 28858
rect 65386 28806 65438 28858
rect 65450 28806 65502 28858
rect 65514 28806 65566 28858
rect 65064 28747 65116 28756
rect 65064 28713 65073 28747
rect 65073 28713 65107 28747
rect 65107 28713 65116 28747
rect 65064 28704 65116 28713
rect 65156 28636 65208 28688
rect 65984 28568 66036 28620
rect 64972 28432 65024 28484
rect 64338 28262 64390 28314
rect 64402 28262 64454 28314
rect 64466 28262 64518 28314
rect 64530 28262 64582 28314
rect 64594 28262 64646 28314
rect 65258 27718 65310 27770
rect 65322 27718 65374 27770
rect 65386 27718 65438 27770
rect 65450 27718 65502 27770
rect 65514 27718 65566 27770
rect 62856 27548 62908 27600
rect 63500 27548 63552 27600
rect 64338 27174 64390 27226
rect 64402 27174 64454 27226
rect 64466 27174 64518 27226
rect 64530 27174 64582 27226
rect 64594 27174 64646 27226
rect 65064 27004 65116 27056
rect 64972 26936 65024 26988
rect 65708 26868 65760 26920
rect 65800 26800 65852 26852
rect 65258 26630 65310 26682
rect 65322 26630 65374 26682
rect 65386 26630 65438 26682
rect 65450 26630 65502 26682
rect 65514 26630 65566 26682
rect 64972 26528 65024 26580
rect 65616 26528 65668 26580
rect 64052 26367 64104 26376
rect 64052 26333 64061 26367
rect 64061 26333 64095 26367
rect 64095 26333 64104 26367
rect 64052 26324 64104 26333
rect 64696 26324 64748 26376
rect 64972 26324 65024 26376
rect 66168 26460 66220 26512
rect 65984 26188 66036 26240
rect 64338 26086 64390 26138
rect 64402 26086 64454 26138
rect 64466 26086 64518 26138
rect 64530 26086 64582 26138
rect 64594 26086 64646 26138
rect 64696 25984 64748 26036
rect 65064 25891 65116 25900
rect 65064 25857 65073 25891
rect 65073 25857 65107 25891
rect 65107 25857 65116 25891
rect 65064 25848 65116 25857
rect 65156 25848 65208 25900
rect 65708 25848 65760 25900
rect 65984 25823 66036 25832
rect 65984 25789 65993 25823
rect 65993 25789 66027 25823
rect 66027 25789 66036 25823
rect 65984 25780 66036 25789
rect 65258 25542 65310 25594
rect 65322 25542 65374 25594
rect 65386 25542 65438 25594
rect 65450 25542 65502 25594
rect 65514 25542 65566 25594
rect 63960 25304 64012 25356
rect 65064 25279 65116 25288
rect 65064 25245 65073 25279
rect 65073 25245 65107 25279
rect 65107 25245 65116 25279
rect 65064 25236 65116 25245
rect 65156 25279 65208 25288
rect 65156 25245 65165 25279
rect 65165 25245 65199 25279
rect 65199 25245 65208 25279
rect 65156 25236 65208 25245
rect 65800 25236 65852 25288
rect 64236 25100 64288 25152
rect 64338 24998 64390 25050
rect 64402 24998 64454 25050
rect 64466 24998 64518 25050
rect 64530 24998 64582 25050
rect 64594 24998 64646 25050
rect 64880 24692 64932 24744
rect 63960 24556 64012 24608
rect 65258 24454 65310 24506
rect 65322 24454 65374 24506
rect 65386 24454 65438 24506
rect 65450 24454 65502 24506
rect 65514 24454 65566 24506
rect 64236 24284 64288 24336
rect 64972 24284 65024 24336
rect 63960 24148 64012 24200
rect 65800 24055 65852 24064
rect 65800 24021 65809 24055
rect 65809 24021 65843 24055
rect 65843 24021 65852 24055
rect 65800 24012 65852 24021
rect 64338 23910 64390 23962
rect 64402 23910 64454 23962
rect 64466 23910 64518 23962
rect 64530 23910 64582 23962
rect 64594 23910 64646 23962
rect 63040 23740 63092 23792
rect 63868 23740 63920 23792
rect 62764 23604 62816 23656
rect 63408 23468 63460 23520
rect 63684 23468 63736 23520
rect 64052 23468 64104 23520
rect 65258 23366 65310 23418
rect 65322 23366 65374 23418
rect 65386 23366 65438 23418
rect 65450 23366 65502 23418
rect 65514 23366 65566 23418
rect 65064 23264 65116 23316
rect 65984 23196 66036 23248
rect 64052 23171 64104 23180
rect 64052 23137 64061 23171
rect 64061 23137 64095 23171
rect 64095 23137 64104 23171
rect 64052 23128 64104 23137
rect 64972 23128 65024 23180
rect 66536 23128 66588 23180
rect 65616 23060 65668 23112
rect 63132 22992 63184 23044
rect 64880 22992 64932 23044
rect 64338 22822 64390 22874
rect 64402 22822 64454 22874
rect 64466 22822 64518 22874
rect 64530 22822 64582 22874
rect 64594 22822 64646 22874
rect 64972 22720 65024 22772
rect 65258 22278 65310 22330
rect 65322 22278 65374 22330
rect 65386 22278 65438 22330
rect 65450 22278 65502 22330
rect 65514 22278 65566 22330
rect 66352 22176 66404 22228
rect 66168 22108 66220 22160
rect 63960 21972 64012 22024
rect 64696 21972 64748 22024
rect 64338 21734 64390 21786
rect 64402 21734 64454 21786
rect 64466 21734 64518 21786
rect 64530 21734 64582 21786
rect 64594 21734 64646 21786
rect 66352 21496 66404 21548
rect 63316 21428 63368 21480
rect 63868 21428 63920 21480
rect 65616 21360 65668 21412
rect 64972 21292 65024 21344
rect 65258 21190 65310 21242
rect 65322 21190 65374 21242
rect 65386 21190 65438 21242
rect 65450 21190 65502 21242
rect 65514 21190 65566 21242
rect 64696 21088 64748 21140
rect 64972 21131 65024 21140
rect 64972 21097 64981 21131
rect 64981 21097 65015 21131
rect 65015 21097 65024 21131
rect 64972 21088 65024 21097
rect 65156 21020 65208 21072
rect 66076 21020 66128 21072
rect 65616 20884 65668 20936
rect 66168 20748 66220 20800
rect 64338 20646 64390 20698
rect 64402 20646 64454 20698
rect 64466 20646 64518 20698
rect 64530 20646 64582 20698
rect 64594 20646 64646 20698
rect 64144 20544 64196 20596
rect 65892 20544 65944 20596
rect 65064 20476 65116 20528
rect 65708 20408 65760 20460
rect 65800 20340 65852 20392
rect 64972 20247 65024 20256
rect 64972 20213 64981 20247
rect 64981 20213 65015 20247
rect 65015 20213 65024 20247
rect 64972 20204 65024 20213
rect 65258 20102 65310 20154
rect 65322 20102 65374 20154
rect 65386 20102 65438 20154
rect 65450 20102 65502 20154
rect 65514 20102 65566 20154
rect 66168 19932 66220 19984
rect 64052 19907 64104 19916
rect 64052 19873 64061 19907
rect 64061 19873 64095 19907
rect 64095 19873 64104 19907
rect 64052 19864 64104 19873
rect 64696 19796 64748 19848
rect 65984 19660 66036 19712
rect 64338 19558 64390 19610
rect 64402 19558 64454 19610
rect 64466 19558 64518 19610
rect 64530 19558 64582 19610
rect 64594 19558 64646 19610
rect 64696 19456 64748 19508
rect 65616 19320 65668 19372
rect 65064 19295 65116 19304
rect 65064 19261 65073 19295
rect 65073 19261 65107 19295
rect 65107 19261 65116 19295
rect 65064 19252 65116 19261
rect 65984 19295 66036 19304
rect 65984 19261 65993 19295
rect 65993 19261 66027 19295
rect 66027 19261 66036 19295
rect 65984 19252 66036 19261
rect 65258 19014 65310 19066
rect 65322 19014 65374 19066
rect 65386 19014 65438 19066
rect 65450 19014 65502 19066
rect 65514 19014 65566 19066
rect 65064 18751 65116 18760
rect 65064 18717 65073 18751
rect 65073 18717 65107 18751
rect 65107 18717 65116 18751
rect 65064 18708 65116 18717
rect 65616 18708 65668 18760
rect 65800 18708 65852 18760
rect 64696 18572 64748 18624
rect 64338 18470 64390 18522
rect 64402 18470 64454 18522
rect 64466 18470 64518 18522
rect 64530 18470 64582 18522
rect 64594 18470 64646 18522
rect 64052 18275 64104 18284
rect 64052 18241 64061 18275
rect 64061 18241 64095 18275
rect 64095 18241 64104 18275
rect 64052 18232 64104 18241
rect 64696 18232 64748 18284
rect 66168 18096 66220 18148
rect 65800 18071 65852 18080
rect 65800 18037 65809 18071
rect 65809 18037 65843 18071
rect 65843 18037 65852 18071
rect 65800 18028 65852 18037
rect 65258 17926 65310 17978
rect 65322 17926 65374 17978
rect 65386 17926 65438 17978
rect 65450 17926 65502 17978
rect 65514 17926 65566 17978
rect 64236 17824 64288 17876
rect 65064 17824 65116 17876
rect 66352 17824 66404 17876
rect 65800 17756 65852 17808
rect 65708 17688 65760 17740
rect 64880 17620 64932 17672
rect 65156 17552 65208 17604
rect 65708 17552 65760 17604
rect 64338 17382 64390 17434
rect 64402 17382 64454 17434
rect 64466 17382 64518 17434
rect 64530 17382 64582 17434
rect 64594 17382 64646 17434
rect 64236 17280 64288 17332
rect 65258 16838 65310 16890
rect 65322 16838 65374 16890
rect 65386 16838 65438 16890
rect 65450 16838 65502 16890
rect 65514 16838 65566 16890
rect 64972 16736 65024 16788
rect 65156 16668 65208 16720
rect 63316 16396 63368 16448
rect 65892 16396 65944 16448
rect 66076 16439 66128 16448
rect 66076 16405 66085 16439
rect 66085 16405 66119 16439
rect 66119 16405 66128 16439
rect 66076 16396 66128 16405
rect 64338 16294 64390 16346
rect 64402 16294 64454 16346
rect 64466 16294 64518 16346
rect 64530 16294 64582 16346
rect 64594 16294 64646 16346
rect 64880 16192 64932 16244
rect 64788 16124 64840 16176
rect 64604 15988 64656 16040
rect 65984 16124 66036 16176
rect 65892 16099 65944 16108
rect 65892 16065 65901 16099
rect 65901 16065 65935 16099
rect 65935 16065 65944 16099
rect 65892 16056 65944 16065
rect 66444 16056 66496 16108
rect 66076 15988 66128 16040
rect 65258 15750 65310 15802
rect 65322 15750 65374 15802
rect 65386 15750 65438 15802
rect 65450 15750 65502 15802
rect 65514 15750 65566 15802
rect 64604 15691 64656 15700
rect 64604 15657 64613 15691
rect 64613 15657 64647 15691
rect 64647 15657 64656 15691
rect 64604 15648 64656 15657
rect 62764 15308 62816 15360
rect 64144 15308 64196 15360
rect 64338 15206 64390 15258
rect 64402 15206 64454 15258
rect 64466 15206 64518 15258
rect 64530 15206 64582 15258
rect 64594 15206 64646 15258
rect 64788 14968 64840 15020
rect 63868 14900 63920 14952
rect 65064 14832 65116 14884
rect 62948 14764 63000 14816
rect 63684 14764 63736 14816
rect 65156 14764 65208 14816
rect 65800 14807 65852 14816
rect 65800 14773 65809 14807
rect 65809 14773 65843 14807
rect 65843 14773 65852 14807
rect 65800 14764 65852 14773
rect 65258 14662 65310 14714
rect 65322 14662 65374 14714
rect 65386 14662 65438 14714
rect 65450 14662 65502 14714
rect 65514 14662 65566 14714
rect 64338 14118 64390 14170
rect 64402 14118 64454 14170
rect 64466 14118 64518 14170
rect 64530 14118 64582 14170
rect 64594 14118 64646 14170
rect 63040 13812 63092 13864
rect 63592 13812 63644 13864
rect 65258 13574 65310 13626
rect 65322 13574 65374 13626
rect 65386 13574 65438 13626
rect 65450 13574 65502 13626
rect 65514 13574 65566 13626
rect 65708 13472 65760 13524
rect 64236 13404 64288 13456
rect 65616 13404 65668 13456
rect 66168 13404 66220 13456
rect 63868 13268 63920 13320
rect 64338 13030 64390 13082
rect 64402 13030 64454 13082
rect 64466 13030 64518 13082
rect 64530 13030 64582 13082
rect 64594 13030 64646 13082
rect 65708 12792 65760 12844
rect 64972 12588 65024 12640
rect 65258 12486 65310 12538
rect 65322 12486 65374 12538
rect 65386 12486 65438 12538
rect 65450 12486 65502 12538
rect 65514 12486 65566 12538
rect 65616 12316 65668 12368
rect 63868 12180 63920 12232
rect 64696 12180 64748 12232
rect 66352 12180 66404 12232
rect 64338 11942 64390 11994
rect 64402 11942 64454 11994
rect 64466 11942 64518 11994
rect 64530 11942 64582 11994
rect 64594 11942 64646 11994
rect 64236 11840 64288 11892
rect 65156 11747 65208 11756
rect 65156 11713 65165 11747
rect 65165 11713 65199 11747
rect 65199 11713 65208 11747
rect 65156 11704 65208 11713
rect 64972 11679 65024 11688
rect 64972 11645 64981 11679
rect 64981 11645 65015 11679
rect 65015 11645 65024 11679
rect 64972 11636 65024 11645
rect 63960 11500 64012 11552
rect 65258 11398 65310 11450
rect 65322 11398 65374 11450
rect 65386 11398 65438 11450
rect 65450 11398 65502 11450
rect 65514 11398 65566 11450
rect 64696 11296 64748 11348
rect 63684 11228 63736 11280
rect 66352 11228 66404 11280
rect 66168 11160 66220 11212
rect 65156 11135 65208 11144
rect 65156 11101 65165 11135
rect 65165 11101 65199 11135
rect 65199 11101 65208 11135
rect 65156 11092 65208 11101
rect 64338 10854 64390 10906
rect 64402 10854 64454 10906
rect 64466 10854 64518 10906
rect 64530 10854 64582 10906
rect 64594 10854 64646 10906
rect 64880 10616 64932 10668
rect 65800 10548 65852 10600
rect 64788 10412 64840 10464
rect 64880 10412 64932 10464
rect 65258 10310 65310 10362
rect 65322 10310 65374 10362
rect 65386 10310 65438 10362
rect 65450 10310 65502 10362
rect 65514 10310 65566 10362
rect 65708 10208 65760 10260
rect 64972 10072 65024 10124
rect 64880 10047 64932 10056
rect 64880 10013 64889 10047
rect 64889 10013 64923 10047
rect 64923 10013 64932 10047
rect 64880 10004 64932 10013
rect 65984 10004 66036 10056
rect 65708 9868 65760 9920
rect 64338 9766 64390 9818
rect 64402 9766 64454 9818
rect 64466 9766 64518 9818
rect 64530 9766 64582 9818
rect 64594 9766 64646 9818
rect 65800 9460 65852 9512
rect 64972 9324 65024 9376
rect 65258 9222 65310 9274
rect 65322 9222 65374 9274
rect 65386 9222 65438 9274
rect 65450 9222 65502 9274
rect 65514 9222 65566 9274
rect 65616 9052 65668 9104
rect 63868 8916 63920 8968
rect 64696 8916 64748 8968
rect 65984 8780 66036 8832
rect 64338 8678 64390 8730
rect 64402 8678 64454 8730
rect 64466 8678 64518 8730
rect 64530 8678 64582 8730
rect 64594 8678 64646 8730
rect 64696 8576 64748 8628
rect 65248 8483 65300 8492
rect 65248 8449 65257 8483
rect 65257 8449 65291 8483
rect 65291 8449 65300 8483
rect 65248 8440 65300 8449
rect 65892 8440 65944 8492
rect 65984 8483 66036 8492
rect 65984 8449 65993 8483
rect 65993 8449 66027 8483
rect 66027 8449 66036 8483
rect 65984 8440 66036 8449
rect 65064 8415 65116 8424
rect 65064 8381 65073 8415
rect 65073 8381 65107 8415
rect 65107 8381 65116 8415
rect 65064 8372 65116 8381
rect 65258 8134 65310 8186
rect 65322 8134 65374 8186
rect 65386 8134 65438 8186
rect 65450 8134 65502 8186
rect 65514 8134 65566 8186
rect 65800 8075 65852 8084
rect 65800 8041 65809 8075
rect 65809 8041 65843 8075
rect 65843 8041 65852 8075
rect 65800 8032 65852 8041
rect 65616 7964 65668 8016
rect 66076 7964 66128 8016
rect 64052 7939 64104 7948
rect 64052 7905 64061 7939
rect 64061 7905 64095 7939
rect 64095 7905 64104 7939
rect 64052 7896 64104 7905
rect 64696 7828 64748 7880
rect 64338 7590 64390 7642
rect 64402 7590 64454 7642
rect 64466 7590 64518 7642
rect 64530 7590 64582 7642
rect 64594 7590 64646 7642
rect 64144 7488 64196 7540
rect 64696 7488 64748 7540
rect 64788 7352 64840 7404
rect 65892 7352 65944 7404
rect 64972 7327 65024 7336
rect 64972 7293 64981 7327
rect 64981 7293 65015 7327
rect 65015 7293 65024 7327
rect 64972 7284 65024 7293
rect 65984 7327 66036 7336
rect 65984 7293 65993 7327
rect 65993 7293 66027 7327
rect 66027 7293 66036 7327
rect 65984 7284 66036 7293
rect 65616 7148 65668 7200
rect 65258 7046 65310 7098
rect 65322 7046 65374 7098
rect 65386 7046 65438 7098
rect 65450 7046 65502 7098
rect 65514 7046 65566 7098
rect 64144 6944 64196 6996
rect 65616 6987 65668 6996
rect 65616 6953 65625 6987
rect 65625 6953 65659 6987
rect 65659 6953 65668 6987
rect 65616 6944 65668 6953
rect 63776 6808 63828 6860
rect 65800 6876 65852 6928
rect 65708 6851 65760 6860
rect 65708 6817 65717 6851
rect 65717 6817 65751 6851
rect 65751 6817 65760 6851
rect 65708 6808 65760 6817
rect 64880 6740 64932 6792
rect 65800 6783 65852 6792
rect 65800 6749 65809 6783
rect 65809 6749 65843 6783
rect 65843 6749 65852 6783
rect 65800 6740 65852 6749
rect 65064 6672 65116 6724
rect 64236 6604 64288 6656
rect 64338 6502 64390 6554
rect 64402 6502 64454 6554
rect 64466 6502 64518 6554
rect 64530 6502 64582 6554
rect 64594 6502 64646 6554
rect 64144 6400 64196 6452
rect 63960 6332 64012 6384
rect 64880 6264 64932 6316
rect 65984 6196 66036 6248
rect 64696 6060 64748 6112
rect 65258 5958 65310 6010
rect 65322 5958 65374 6010
rect 65386 5958 65438 6010
rect 65450 5958 65502 6010
rect 65514 5958 65566 6010
rect 64144 5899 64196 5908
rect 64144 5865 64153 5899
rect 64153 5865 64187 5899
rect 64187 5865 64196 5899
rect 64144 5856 64196 5865
rect 64696 5899 64748 5908
rect 64696 5865 64705 5899
rect 64705 5865 64739 5899
rect 64739 5865 64748 5899
rect 64696 5856 64748 5865
rect 64880 5856 64932 5908
rect 65432 5856 65484 5908
rect 65800 5856 65852 5908
rect 65708 5788 65760 5840
rect 63960 5652 64012 5704
rect 64788 5720 64840 5772
rect 65064 5720 65116 5772
rect 64696 5652 64748 5704
rect 65432 5695 65484 5704
rect 65432 5661 65441 5695
rect 65441 5661 65475 5695
rect 65475 5661 65484 5695
rect 65432 5652 65484 5661
rect 64972 5584 65024 5636
rect 64788 5516 64840 5568
rect 64338 5414 64390 5466
rect 64402 5414 64454 5466
rect 64466 5414 64518 5466
rect 64530 5414 64582 5466
rect 64594 5414 64646 5466
rect 63868 5219 63920 5228
rect 63868 5185 63877 5219
rect 63877 5185 63911 5219
rect 63911 5185 63920 5219
rect 63868 5176 63920 5185
rect 64788 5176 64840 5228
rect 65616 5108 65668 5160
rect 66076 5108 66128 5160
rect 65708 4972 65760 5024
rect 65258 4870 65310 4922
rect 65322 4870 65374 4922
rect 65386 4870 65438 4922
rect 65450 4870 65502 4922
rect 65514 4870 65566 4922
rect 65984 4768 66036 4820
rect 64236 4700 64288 4752
rect 65616 4700 65668 4752
rect 64052 4675 64104 4684
rect 64052 4641 64061 4675
rect 64061 4641 64095 4675
rect 64095 4641 64104 4675
rect 64052 4632 64104 4641
rect 64338 4326 64390 4378
rect 64402 4326 64454 4378
rect 64466 4326 64518 4378
rect 64530 4326 64582 4378
rect 64594 4326 64646 4378
rect 63408 4224 63460 4276
rect 64236 4224 64288 4276
rect 64052 3952 64104 4004
rect 64144 3995 64196 4004
rect 64144 3961 64153 3995
rect 64153 3961 64187 3995
rect 64187 3961 64196 3995
rect 64144 3952 64196 3961
rect 65156 3952 65208 4004
rect 65984 3884 66036 3936
rect 65258 3782 65310 3834
rect 65322 3782 65374 3834
rect 65386 3782 65438 3834
rect 65450 3782 65502 3834
rect 65514 3782 65566 3834
rect 64144 3680 64196 3732
rect 64236 3655 64288 3664
rect 64236 3621 64245 3655
rect 64245 3621 64279 3655
rect 64279 3621 64288 3655
rect 64236 3612 64288 3621
rect 65156 3612 65208 3664
rect 63960 3519 64012 3528
rect 63960 3485 63969 3519
rect 63969 3485 64003 3519
rect 64003 3485 64012 3519
rect 63960 3476 64012 3485
rect 64696 3408 64748 3460
rect 64972 3476 65024 3528
rect 66444 3476 66496 3528
rect 65984 3408 66036 3460
rect 63776 3340 63828 3392
rect 64788 3340 64840 3392
rect 64338 3238 64390 3290
rect 64402 3238 64454 3290
rect 64466 3238 64518 3290
rect 64530 3238 64582 3290
rect 64594 3238 64646 3290
rect 64144 3136 64196 3188
rect 64052 3043 64104 3052
rect 64052 3009 64061 3043
rect 64061 3009 64095 3043
rect 64095 3009 64104 3043
rect 64052 3000 64104 3009
rect 65800 3043 65852 3052
rect 65800 3009 65809 3043
rect 65809 3009 65843 3043
rect 65843 3009 65852 3043
rect 65800 3000 65852 3009
rect 64328 2907 64380 2916
rect 64328 2873 64337 2907
rect 64337 2873 64371 2907
rect 64371 2873 64380 2907
rect 64328 2864 64380 2873
rect 65616 2864 65668 2916
rect 65258 2694 65310 2746
rect 65322 2694 65374 2746
rect 65386 2694 65438 2746
rect 65450 2694 65502 2746
rect 65514 2694 65566 2746
rect 64328 2592 64380 2644
rect 65708 2592 65760 2644
rect 66352 2524 66404 2576
rect 64972 2456 65024 2508
rect 64788 2388 64840 2440
rect 65248 2431 65300 2440
rect 65248 2397 65257 2431
rect 65257 2397 65291 2431
rect 65291 2397 65300 2431
rect 65248 2388 65300 2397
rect 64880 2252 64932 2304
rect 64338 2150 64390 2202
rect 64402 2150 64454 2202
rect 64466 2150 64518 2202
rect 64530 2150 64582 2202
rect 64594 2150 64646 2202
rect 65064 2048 65116 2100
rect 49240 1980 49292 2032
rect 62764 1980 62816 2032
rect 66168 1980 66220 2032
rect 48964 1912 49016 1964
rect 62672 1912 62724 1964
rect 65248 1955 65300 1964
rect 65248 1921 65257 1955
rect 65257 1921 65291 1955
rect 65291 1921 65300 1955
rect 65248 1912 65300 1921
rect 65708 1912 65760 1964
rect 49700 1844 49752 1896
rect 63040 1844 63092 1896
rect 64696 1844 64748 1896
rect 65800 1844 65852 1896
rect 65258 1606 65310 1658
rect 65322 1606 65374 1658
rect 65386 1606 65438 1658
rect 65450 1606 65502 1658
rect 65514 1606 65566 1658
rect 65156 1504 65208 1556
rect 64696 1343 64748 1352
rect 64696 1309 64705 1343
rect 64705 1309 64739 1343
rect 64739 1309 64748 1343
rect 64696 1300 64748 1309
rect 65984 1343 66036 1352
rect 65984 1309 65993 1343
rect 65993 1309 66027 1343
rect 66027 1309 66036 1343
rect 65984 1300 66036 1309
rect 64338 1062 64390 1114
rect 64402 1062 64454 1114
rect 64466 1062 64518 1114
rect 64530 1062 64582 1114
rect 64594 1062 64646 1114
rect 64972 960 65024 1012
rect 65800 824 65852 876
rect 65258 518 65310 570
rect 65322 518 65374 570
rect 65386 518 65438 570
rect 65450 518 65502 570
rect 65514 518 65566 570
<< metal2 >>
rect 35346 45112 35402 45121
rect 35346 45047 35402 45056
rect 24858 44976 24914 44985
rect 24858 44911 24914 44920
rect 24872 44810 24900 44911
rect 27712 44872 27764 44878
rect 27712 44814 27764 44820
rect 28816 44872 28868 44878
rect 28816 44814 28868 44820
rect 30932 44872 30984 44878
rect 30932 44814 30984 44820
rect 31758 44840 31814 44849
rect 16764 44804 16816 44810
rect 16764 44746 16816 44752
rect 21732 44804 21784 44810
rect 21732 44746 21784 44752
rect 24860 44804 24912 44810
rect 24860 44746 24912 44752
rect 12530 44704 12586 44713
rect 1998 44636 2306 44645
rect 12530 44639 12586 44648
rect 16210 44704 16266 44713
rect 16210 44639 16266 44648
rect 1998 44634 2004 44636
rect 2060 44634 2084 44636
rect 2140 44634 2164 44636
rect 2220 44634 2244 44636
rect 2300 44634 2306 44636
rect 2060 44582 2062 44634
rect 2242 44582 2244 44634
rect 1998 44580 2004 44582
rect 2060 44580 2084 44582
rect 2140 44580 2164 44582
rect 2220 44580 2244 44582
rect 2300 44580 2306 44582
rect 1998 44571 2306 44580
rect 6182 44568 6238 44577
rect 6182 44503 6184 44512
rect 6236 44503 6238 44512
rect 6734 44568 6790 44577
rect 6734 44503 6736 44512
rect 6184 44474 6236 44480
rect 6788 44503 6790 44512
rect 7286 44568 7342 44577
rect 7286 44503 7288 44512
rect 6736 44474 6788 44480
rect 7340 44503 7342 44512
rect 7838 44568 7894 44577
rect 7838 44503 7840 44512
rect 7288 44474 7340 44480
rect 7892 44503 7894 44512
rect 8390 44568 8446 44577
rect 8390 44503 8392 44512
rect 7840 44474 7892 44480
rect 8444 44503 8446 44512
rect 8942 44568 8998 44577
rect 8942 44503 8944 44512
rect 8392 44474 8444 44480
rect 8996 44503 8998 44512
rect 9494 44568 9550 44577
rect 9494 44503 9496 44512
rect 8944 44474 8996 44480
rect 9548 44503 9550 44512
rect 10046 44568 10102 44577
rect 10046 44503 10048 44512
rect 9496 44474 9548 44480
rect 10100 44503 10102 44512
rect 10598 44568 10654 44577
rect 10598 44503 10600 44512
rect 10048 44474 10100 44480
rect 10652 44503 10654 44512
rect 12254 44568 12310 44577
rect 12544 44538 12572 44639
rect 12806 44568 12862 44577
rect 12254 44503 12256 44512
rect 10600 44474 10652 44480
rect 12308 44503 12310 44512
rect 12532 44532 12584 44538
rect 12256 44474 12308 44480
rect 12806 44503 12808 44512
rect 12532 44474 12584 44480
rect 12860 44503 12862 44512
rect 13542 44568 13598 44577
rect 13542 44503 13544 44512
rect 12808 44474 12860 44480
rect 13596 44503 13598 44512
rect 13818 44568 13874 44577
rect 13818 44503 13820 44512
rect 13544 44474 13596 44480
rect 13872 44503 13874 44512
rect 15474 44568 15530 44577
rect 15474 44503 15476 44512
rect 13820 44474 13872 44480
rect 15528 44503 15530 44512
rect 15934 44568 15990 44577
rect 16224 44538 16252 44639
rect 16670 44568 16726 44577
rect 15934 44503 15936 44512
rect 15476 44474 15528 44480
rect 15988 44503 15990 44512
rect 16212 44532 16264 44538
rect 15936 44474 15988 44480
rect 16670 44503 16672 44512
rect 16212 44474 16264 44480
rect 16724 44503 16726 44512
rect 16672 44474 16724 44480
rect 16776 44418 16804 44746
rect 17316 44736 17368 44742
rect 17222 44704 17278 44713
rect 17316 44678 17368 44684
rect 17222 44639 17278 44648
rect 16946 44568 17002 44577
rect 17236 44538 17264 44639
rect 16946 44503 16948 44512
rect 17000 44503 17002 44512
rect 17224 44532 17276 44538
rect 16948 44474 17000 44480
rect 17224 44474 17276 44480
rect 16684 44390 16804 44418
rect 12256 44328 12308 44334
rect 12256 44270 12308 44276
rect 14372 44328 14424 44334
rect 14372 44270 14424 44276
rect 10600 44260 10652 44266
rect 10600 44202 10652 44208
rect 2918 44092 3226 44101
rect 2918 44090 2924 44092
rect 2980 44090 3004 44092
rect 3060 44090 3084 44092
rect 3140 44090 3164 44092
rect 3220 44090 3226 44092
rect 2980 44038 2982 44090
rect 3162 44038 3164 44090
rect 2918 44036 2924 44038
rect 2980 44036 3004 44038
rect 3060 44036 3084 44038
rect 3140 44036 3164 44038
rect 3220 44036 3226 44038
rect 2918 44027 3226 44036
rect 1998 43548 2306 43557
rect 1998 43546 2004 43548
rect 2060 43546 2084 43548
rect 2140 43546 2164 43548
rect 2220 43546 2244 43548
rect 2300 43546 2306 43548
rect 2060 43494 2062 43546
rect 2242 43494 2244 43546
rect 1998 43492 2004 43494
rect 2060 43492 2084 43494
rect 2140 43492 2164 43494
rect 2220 43492 2244 43494
rect 2300 43492 2306 43494
rect 1998 43483 2306 43492
rect 10612 43178 10640 44202
rect 11612 44192 11664 44198
rect 11612 44134 11664 44140
rect 11624 43994 11652 44134
rect 11612 43988 11664 43994
rect 11612 43930 11664 43936
rect 11150 43888 11206 43897
rect 11150 43823 11152 43832
rect 11204 43823 11206 43832
rect 11152 43794 11204 43800
rect 11060 43648 11112 43654
rect 11060 43590 11112 43596
rect 11072 43314 11100 43590
rect 11060 43308 11112 43314
rect 11060 43250 11112 43256
rect 10600 43172 10652 43178
rect 10600 43114 10652 43120
rect 11704 43172 11756 43178
rect 11704 43114 11756 43120
rect 2918 43004 3226 43013
rect 2918 43002 2924 43004
rect 2980 43002 3004 43004
rect 3060 43002 3084 43004
rect 3140 43002 3164 43004
rect 3220 43002 3226 43004
rect 2980 42950 2982 43002
rect 3162 42950 3164 43002
rect 2918 42948 2924 42950
rect 2980 42948 3004 42950
rect 3060 42948 3084 42950
rect 3140 42948 3164 42950
rect 3220 42948 3226 42950
rect 2918 42939 3226 42948
rect 1998 42460 2306 42469
rect 1998 42458 2004 42460
rect 2060 42458 2084 42460
rect 2140 42458 2164 42460
rect 2220 42458 2244 42460
rect 2300 42458 2306 42460
rect 2060 42406 2062 42458
rect 2242 42406 2244 42458
rect 1998 42404 2004 42406
rect 2060 42404 2084 42406
rect 2140 42404 2164 42406
rect 2220 42404 2244 42406
rect 2300 42404 2306 42406
rect 1998 42395 2306 42404
rect 10416 42356 10468 42362
rect 10416 42298 10468 42304
rect 7932 42152 7984 42158
rect 7932 42094 7984 42100
rect 9772 42152 9824 42158
rect 9772 42094 9824 42100
rect 2918 41916 3226 41925
rect 2918 41914 2924 41916
rect 2980 41914 3004 41916
rect 3060 41914 3084 41916
rect 3140 41914 3164 41916
rect 3220 41914 3226 41916
rect 2980 41862 2982 41914
rect 3162 41862 3164 41914
rect 2918 41860 2924 41862
rect 2980 41860 3004 41862
rect 3060 41860 3084 41862
rect 3140 41860 3164 41862
rect 3220 41860 3226 41862
rect 2918 41851 3226 41860
rect 7944 41614 7972 42094
rect 9784 41750 9812 42094
rect 10428 41818 10456 42298
rect 10612 42226 10640 43114
rect 11716 42906 11744 43114
rect 12268 43092 12296 44270
rect 14188 44260 14240 44266
rect 14188 44202 14240 44208
rect 12532 44192 12584 44198
rect 12452 44152 12532 44180
rect 12452 43790 12480 44152
rect 12532 44134 12584 44140
rect 12900 44192 12952 44198
rect 12900 44134 12952 44140
rect 12532 43852 12584 43858
rect 12532 43794 12584 43800
rect 12440 43784 12492 43790
rect 12440 43726 12492 43732
rect 12348 43104 12400 43110
rect 12268 43064 12348 43092
rect 12268 42906 12296 43064
rect 12348 43046 12400 43052
rect 12544 42906 12572 43794
rect 12716 43648 12768 43654
rect 12716 43590 12768 43596
rect 12728 43450 12756 43590
rect 12716 43444 12768 43450
rect 12716 43386 12768 43392
rect 11704 42900 11756 42906
rect 11704 42842 11756 42848
rect 12256 42900 12308 42906
rect 12256 42842 12308 42848
rect 12532 42900 12584 42906
rect 12532 42842 12584 42848
rect 10600 42220 10652 42226
rect 10600 42162 10652 42168
rect 10968 42220 11020 42226
rect 10968 42162 11020 42168
rect 10692 42016 10744 42022
rect 10692 41958 10744 41964
rect 10416 41812 10468 41818
rect 10416 41754 10468 41760
rect 9772 41744 9824 41750
rect 9772 41686 9824 41692
rect 7932 41608 7984 41614
rect 7932 41550 7984 41556
rect 8208 41608 8260 41614
rect 8208 41550 8260 41556
rect 1998 41372 2306 41381
rect 1998 41370 2004 41372
rect 2060 41370 2084 41372
rect 2140 41370 2164 41372
rect 2220 41370 2244 41372
rect 2300 41370 2306 41372
rect 2060 41318 2062 41370
rect 2242 41318 2244 41370
rect 1998 41316 2004 41318
rect 2060 41316 2084 41318
rect 2140 41316 2164 41318
rect 2220 41316 2244 41318
rect 2300 41316 2306 41318
rect 1998 41307 2306 41316
rect 2918 40828 3226 40837
rect 2918 40826 2924 40828
rect 2980 40826 3004 40828
rect 3060 40826 3084 40828
rect 3140 40826 3164 40828
rect 3220 40826 3226 40828
rect 2980 40774 2982 40826
rect 3162 40774 3164 40826
rect 2918 40772 2924 40774
rect 2980 40772 3004 40774
rect 3060 40772 3084 40774
rect 3140 40772 3164 40774
rect 3220 40772 3226 40774
rect 2918 40763 3226 40772
rect 1998 40284 2306 40293
rect 1998 40282 2004 40284
rect 2060 40282 2084 40284
rect 2140 40282 2164 40284
rect 2220 40282 2244 40284
rect 2300 40282 2306 40284
rect 2060 40230 2062 40282
rect 2242 40230 2244 40282
rect 1998 40228 2004 40230
rect 2060 40228 2084 40230
rect 2140 40228 2164 40230
rect 2220 40228 2244 40230
rect 2300 40228 2306 40230
rect 1998 40219 2306 40228
rect 7944 39982 7972 41550
rect 7932 39976 7984 39982
rect 7932 39918 7984 39924
rect 2918 39740 3226 39749
rect 2918 39738 2924 39740
rect 2980 39738 3004 39740
rect 3060 39738 3084 39740
rect 3140 39738 3164 39740
rect 3220 39738 3226 39740
rect 2980 39686 2982 39738
rect 3162 39686 3164 39738
rect 2918 39684 2924 39686
rect 2980 39684 3004 39686
rect 3060 39684 3084 39686
rect 3140 39684 3164 39686
rect 3220 39684 3226 39686
rect 2918 39675 3226 39684
rect 7840 39296 7892 39302
rect 7840 39238 7892 39244
rect 1998 39196 2306 39205
rect 1998 39194 2004 39196
rect 2060 39194 2084 39196
rect 2140 39194 2164 39196
rect 2220 39194 2244 39196
rect 2300 39194 2306 39196
rect 2060 39142 2062 39194
rect 2242 39142 2244 39194
rect 1998 39140 2004 39142
rect 2060 39140 2084 39142
rect 2140 39140 2164 39142
rect 2220 39140 2244 39142
rect 2300 39140 2306 39142
rect 1998 39131 2306 39140
rect 7104 38956 7156 38962
rect 7104 38898 7156 38904
rect 6920 38752 6972 38758
rect 6920 38694 6972 38700
rect 7012 38752 7064 38758
rect 7012 38694 7064 38700
rect 2918 38652 3226 38661
rect 2918 38650 2924 38652
rect 2980 38650 3004 38652
rect 3060 38650 3084 38652
rect 3140 38650 3164 38652
rect 3220 38650 3226 38652
rect 2980 38598 2982 38650
rect 3162 38598 3164 38650
rect 2918 38596 2924 38598
rect 2980 38596 3004 38598
rect 3060 38596 3084 38598
rect 3140 38596 3164 38598
rect 3220 38596 3226 38598
rect 2918 38587 3226 38596
rect 6932 38554 6960 38694
rect 6920 38548 6972 38554
rect 6920 38490 6972 38496
rect 1998 38108 2306 38117
rect 1998 38106 2004 38108
rect 2060 38106 2084 38108
rect 2140 38106 2164 38108
rect 2220 38106 2244 38108
rect 2300 38106 2306 38108
rect 2060 38054 2062 38106
rect 2242 38054 2244 38106
rect 1998 38052 2004 38054
rect 2060 38052 2084 38054
rect 2140 38052 2164 38054
rect 2220 38052 2244 38054
rect 2300 38052 2306 38054
rect 1998 38043 2306 38052
rect 7024 37738 7052 38694
rect 7116 37874 7144 38898
rect 7852 38554 7880 39238
rect 7944 38962 7972 39918
rect 8220 39846 8248 41550
rect 9680 41472 9732 41478
rect 9680 41414 9732 41420
rect 8760 41132 8812 41138
rect 8760 41074 8812 41080
rect 8772 40526 8800 41074
rect 9692 41002 9720 41414
rect 9784 41002 9812 41686
rect 10416 41608 10468 41614
rect 10416 41550 10468 41556
rect 10048 41472 10100 41478
rect 10048 41414 10100 41420
rect 10060 41138 10088 41414
rect 10048 41132 10100 41138
rect 10048 41074 10100 41080
rect 9680 40996 9732 41002
rect 9680 40938 9732 40944
rect 9772 40996 9824 41002
rect 9772 40938 9824 40944
rect 10140 40996 10192 41002
rect 10140 40938 10192 40944
rect 8944 40928 8996 40934
rect 8944 40870 8996 40876
rect 8760 40520 8812 40526
rect 8760 40462 8812 40468
rect 8208 39840 8260 39846
rect 8208 39782 8260 39788
rect 8208 39432 8260 39438
rect 8208 39374 8260 39380
rect 8220 39098 8248 39374
rect 8208 39092 8260 39098
rect 8208 39034 8260 39040
rect 7932 38956 7984 38962
rect 7932 38898 7984 38904
rect 8220 38554 8248 39034
rect 8392 38956 8444 38962
rect 8392 38898 8444 38904
rect 7840 38548 7892 38554
rect 7840 38490 7892 38496
rect 8208 38548 8260 38554
rect 8208 38490 8260 38496
rect 8404 38418 8432 38898
rect 8772 38554 8800 40462
rect 8956 39914 8984 40870
rect 9036 40520 9088 40526
rect 9036 40462 9088 40468
rect 9048 40186 9076 40462
rect 9036 40180 9088 40186
rect 9036 40122 9088 40128
rect 9312 40044 9364 40050
rect 9312 39986 9364 39992
rect 8944 39908 8996 39914
rect 8944 39850 8996 39856
rect 9324 38962 9352 39986
rect 9692 39846 9720 40938
rect 10152 40594 10180 40938
rect 10140 40588 10192 40594
rect 10140 40530 10192 40536
rect 10324 40588 10376 40594
rect 10324 40530 10376 40536
rect 9772 40520 9824 40526
rect 9772 40462 9824 40468
rect 9680 39840 9732 39846
rect 9680 39782 9732 39788
rect 9784 39658 9812 40462
rect 10336 40118 10364 40530
rect 10324 40112 10376 40118
rect 10324 40054 10376 40060
rect 10428 40050 10456 41550
rect 10704 40730 10732 41958
rect 10980 41546 11008 42162
rect 11428 41676 11480 41682
rect 11428 41618 11480 41624
rect 11336 41608 11388 41614
rect 11336 41550 11388 41556
rect 10968 41540 11020 41546
rect 10968 41482 11020 41488
rect 10784 41472 10836 41478
rect 10784 41414 10836 41420
rect 10692 40724 10744 40730
rect 10692 40666 10744 40672
rect 10416 40044 10468 40050
rect 10416 39986 10468 39992
rect 10140 39840 10192 39846
rect 10140 39782 10192 39788
rect 9692 39630 9812 39658
rect 9692 39574 9720 39630
rect 10152 39574 10180 39782
rect 9680 39568 9732 39574
rect 9680 39510 9732 39516
rect 10140 39568 10192 39574
rect 10140 39510 10192 39516
rect 9312 38956 9364 38962
rect 9312 38898 9364 38904
rect 9692 38894 9720 39510
rect 10428 39370 10456 39986
rect 10692 39840 10744 39846
rect 10796 39828 10824 41414
rect 10980 40186 11008 41482
rect 10968 40180 11020 40186
rect 10968 40122 11020 40128
rect 10744 39800 10824 39828
rect 11060 39840 11112 39846
rect 10692 39782 10744 39788
rect 11060 39782 11112 39788
rect 10416 39364 10468 39370
rect 10416 39306 10468 39312
rect 10324 39296 10376 39302
rect 10324 39238 10376 39244
rect 10336 38962 10364 39238
rect 10324 38956 10376 38962
rect 10324 38898 10376 38904
rect 9680 38888 9732 38894
rect 9680 38830 9732 38836
rect 9956 38888 10008 38894
rect 9956 38830 10008 38836
rect 9864 38752 9916 38758
rect 9864 38694 9916 38700
rect 8760 38548 8812 38554
rect 8760 38490 8812 38496
rect 8392 38412 8444 38418
rect 8392 38354 8444 38360
rect 8484 38412 8536 38418
rect 8484 38354 8536 38360
rect 7380 38344 7432 38350
rect 7380 38286 7432 38292
rect 7932 38344 7984 38350
rect 7932 38286 7984 38292
rect 7392 38010 7420 38286
rect 7380 38004 7432 38010
rect 7380 37946 7432 37952
rect 7944 37942 7972 38286
rect 7932 37936 7984 37942
rect 7932 37878 7984 37884
rect 7104 37868 7156 37874
rect 7104 37810 7156 37816
rect 7012 37732 7064 37738
rect 7012 37674 7064 37680
rect 2918 37564 3226 37573
rect 2918 37562 2924 37564
rect 2980 37562 3004 37564
rect 3060 37562 3084 37564
rect 3140 37562 3164 37564
rect 3220 37562 3226 37564
rect 2980 37510 2982 37562
rect 3162 37510 3164 37562
rect 2918 37508 2924 37510
rect 2980 37508 3004 37510
rect 3060 37508 3084 37510
rect 3140 37508 3164 37510
rect 3220 37508 3226 37510
rect 2918 37499 3226 37508
rect 8496 37330 8524 38354
rect 9876 38010 9904 38694
rect 9968 38418 9996 38830
rect 10232 38820 10284 38826
rect 10232 38762 10284 38768
rect 10324 38820 10376 38826
rect 10324 38762 10376 38768
rect 10244 38486 10272 38762
rect 10232 38480 10284 38486
rect 10232 38422 10284 38428
rect 10336 38418 10364 38762
rect 10968 38752 11020 38758
rect 10968 38694 11020 38700
rect 10980 38554 11008 38694
rect 11072 38554 11100 39782
rect 11348 39506 11376 41550
rect 11440 41138 11468 41618
rect 12912 41614 12940 44134
rect 12992 43920 13044 43926
rect 12992 43862 13044 43868
rect 13004 43178 13032 43862
rect 14004 43444 14056 43450
rect 14004 43386 14056 43392
rect 12992 43172 13044 43178
rect 12992 43114 13044 43120
rect 13820 43172 13872 43178
rect 13820 43114 13872 43120
rect 12624 41608 12676 41614
rect 12624 41550 12676 41556
rect 12900 41608 12952 41614
rect 12900 41550 12952 41556
rect 11888 41472 11940 41478
rect 11888 41414 11940 41420
rect 11428 41132 11480 41138
rect 11428 41074 11480 41080
rect 11440 40934 11468 41074
rect 11900 41002 11928 41414
rect 12440 41132 12492 41138
rect 12440 41074 12492 41080
rect 11888 40996 11940 41002
rect 11888 40938 11940 40944
rect 11428 40928 11480 40934
rect 11428 40870 11480 40876
rect 11440 40730 11468 40870
rect 11428 40724 11480 40730
rect 11428 40666 11480 40672
rect 11426 40624 11482 40633
rect 11426 40559 11428 40568
rect 11480 40559 11482 40568
rect 11428 40530 11480 40536
rect 11440 39914 11468 40530
rect 12256 40520 12308 40526
rect 12256 40462 12308 40468
rect 11428 39908 11480 39914
rect 11428 39850 11480 39856
rect 11612 39840 11664 39846
rect 11612 39782 11664 39788
rect 11624 39681 11652 39782
rect 11610 39672 11666 39681
rect 11440 39630 11610 39658
rect 11336 39500 11388 39506
rect 11336 39442 11388 39448
rect 10968 38548 11020 38554
rect 10968 38490 11020 38496
rect 11060 38548 11112 38554
rect 11060 38490 11112 38496
rect 11440 38418 11468 39630
rect 11610 39607 11666 39616
rect 12072 39500 12124 39506
rect 12072 39442 12124 39448
rect 11612 39432 11664 39438
rect 11612 39374 11664 39380
rect 9956 38412 10008 38418
rect 9956 38354 10008 38360
rect 10324 38412 10376 38418
rect 10324 38354 10376 38360
rect 11428 38412 11480 38418
rect 11428 38354 11480 38360
rect 11520 38344 11572 38350
rect 11520 38286 11572 38292
rect 9956 38276 10008 38282
rect 9956 38218 10008 38224
rect 9864 38004 9916 38010
rect 9864 37946 9916 37952
rect 9036 37732 9088 37738
rect 9036 37674 9088 37680
rect 8760 37664 8812 37670
rect 8760 37606 8812 37612
rect 8772 37398 8800 37606
rect 9048 37398 9076 37674
rect 9968 37670 9996 38218
rect 11532 37806 11560 38286
rect 11624 38282 11652 39374
rect 12084 38826 12112 39442
rect 12268 39030 12296 40462
rect 12452 39982 12480 41074
rect 12440 39976 12492 39982
rect 12440 39918 12492 39924
rect 12452 39302 12480 39918
rect 12636 39846 12664 41550
rect 13004 41414 13032 43114
rect 13176 43104 13228 43110
rect 13176 43046 13228 43052
rect 13188 42770 13216 43046
rect 13176 42764 13228 42770
rect 13176 42706 13228 42712
rect 13084 42696 13136 42702
rect 13084 42638 13136 42644
rect 13544 42696 13596 42702
rect 13544 42638 13596 42644
rect 12912 41386 13032 41414
rect 12912 41002 12940 41386
rect 13096 41206 13124 42638
rect 13556 42362 13584 42638
rect 13832 42634 13860 43114
rect 14016 42906 14044 43386
rect 14004 42900 14056 42906
rect 14004 42842 14056 42848
rect 14016 42702 14044 42842
rect 14200 42838 14228 44202
rect 14384 43994 14412 44270
rect 14740 44192 14792 44198
rect 14740 44134 14792 44140
rect 14832 44192 14884 44198
rect 14832 44134 14884 44140
rect 14372 43988 14424 43994
rect 14372 43930 14424 43936
rect 14280 43172 14332 43178
rect 14280 43114 14332 43120
rect 14188 42832 14240 42838
rect 14188 42774 14240 42780
rect 14004 42696 14056 42702
rect 14004 42638 14056 42644
rect 13820 42628 13872 42634
rect 13820 42570 13872 42576
rect 14200 42378 14228 42774
rect 14292 42566 14320 43114
rect 14384 42906 14412 43930
rect 14752 43858 14780 44134
rect 14844 43994 14872 44134
rect 14832 43988 14884 43994
rect 14832 43930 14884 43936
rect 16120 43988 16172 43994
rect 16120 43930 16172 43936
rect 15290 43888 15346 43897
rect 14740 43852 14792 43858
rect 15290 43823 15292 43832
rect 14740 43794 14792 43800
rect 15344 43823 15346 43832
rect 15660 43852 15712 43858
rect 15292 43794 15344 43800
rect 15660 43794 15712 43800
rect 14740 43648 14792 43654
rect 14740 43590 14792 43596
rect 14752 42906 14780 43590
rect 15568 43104 15620 43110
rect 15568 43046 15620 43052
rect 14372 42900 14424 42906
rect 14372 42842 14424 42848
rect 14740 42900 14792 42906
rect 14740 42842 14792 42848
rect 14556 42764 14608 42770
rect 14556 42706 14608 42712
rect 14280 42560 14332 42566
rect 14280 42502 14332 42508
rect 13544 42356 13596 42362
rect 14200 42350 14320 42378
rect 13544 42298 13596 42304
rect 14188 42220 14240 42226
rect 14188 42162 14240 42168
rect 13820 41608 13872 41614
rect 13820 41550 13872 41556
rect 13176 41540 13228 41546
rect 13176 41482 13228 41488
rect 13084 41200 13136 41206
rect 13084 41142 13136 41148
rect 12900 40996 12952 41002
rect 12900 40938 12952 40944
rect 12808 40928 12860 40934
rect 12808 40870 12860 40876
rect 12820 40050 12848 40870
rect 12808 40044 12860 40050
rect 12808 39986 12860 39992
rect 12714 39944 12770 39953
rect 12714 39879 12770 39888
rect 12624 39840 12676 39846
rect 12624 39782 12676 39788
rect 12532 39432 12584 39438
rect 12532 39374 12584 39380
rect 12440 39296 12492 39302
rect 12440 39238 12492 39244
rect 12544 39098 12572 39374
rect 12532 39092 12584 39098
rect 12532 39034 12584 39040
rect 12256 39024 12308 39030
rect 12256 38966 12308 38972
rect 12072 38820 12124 38826
rect 12072 38762 12124 38768
rect 12084 38457 12112 38762
rect 12070 38448 12126 38457
rect 12070 38383 12072 38392
rect 12124 38383 12126 38392
rect 12072 38354 12124 38360
rect 11612 38276 11664 38282
rect 11612 38218 11664 38224
rect 11520 37800 11572 37806
rect 11520 37742 11572 37748
rect 12084 37738 12112 38354
rect 12268 38350 12296 38966
rect 12728 38418 12756 39879
rect 12912 39574 12940 40938
rect 12900 39568 12952 39574
rect 12900 39510 12952 39516
rect 13188 38962 13216 41482
rect 13728 41268 13780 41274
rect 13728 41210 13780 41216
rect 13740 40916 13768 41210
rect 13832 41070 13860 41550
rect 13820 41064 13872 41070
rect 13820 41006 13872 41012
rect 13820 40928 13872 40934
rect 13740 40888 13820 40916
rect 13740 40526 13768 40888
rect 13820 40870 13872 40876
rect 14096 40928 14148 40934
rect 14096 40870 14148 40876
rect 14108 40662 14136 40870
rect 14096 40656 14148 40662
rect 14096 40598 14148 40604
rect 13728 40520 13780 40526
rect 13728 40462 13780 40468
rect 13740 39982 13768 40462
rect 14200 40050 14228 42162
rect 14188 40044 14240 40050
rect 14188 39986 14240 39992
rect 13728 39976 13780 39982
rect 13728 39918 13780 39924
rect 14200 39642 14228 39986
rect 14188 39636 14240 39642
rect 14188 39578 14240 39584
rect 13820 39364 13872 39370
rect 13820 39306 13872 39312
rect 13544 39296 13596 39302
rect 13544 39238 13596 39244
rect 13176 38956 13228 38962
rect 13176 38898 13228 38904
rect 12716 38412 12768 38418
rect 12716 38354 12768 38360
rect 12164 38344 12216 38350
rect 12164 38286 12216 38292
rect 12256 38344 12308 38350
rect 12256 38286 12308 38292
rect 12808 38344 12860 38350
rect 12808 38286 12860 38292
rect 12072 37732 12124 37738
rect 12072 37674 12124 37680
rect 9956 37664 10008 37670
rect 9956 37606 10008 37612
rect 10508 37664 10560 37670
rect 10508 37606 10560 37612
rect 8760 37392 8812 37398
rect 8760 37334 8812 37340
rect 9036 37392 9088 37398
rect 9036 37334 9088 37340
rect 10520 37330 10548 37606
rect 8484 37324 8536 37330
rect 8484 37266 8536 37272
rect 10508 37324 10560 37330
rect 10508 37266 10560 37272
rect 1998 37020 2306 37029
rect 1998 37018 2004 37020
rect 2060 37018 2084 37020
rect 2140 37018 2164 37020
rect 2220 37018 2244 37020
rect 2300 37018 2306 37020
rect 2060 36966 2062 37018
rect 2242 36966 2244 37018
rect 1998 36964 2004 36966
rect 2060 36964 2084 36966
rect 2140 36964 2164 36966
rect 2220 36964 2244 36966
rect 2300 36964 2306 36966
rect 1998 36955 2306 36964
rect 10520 36922 10548 37266
rect 10508 36916 10560 36922
rect 10508 36858 10560 36864
rect 12176 36009 12204 38286
rect 12268 37874 12296 38286
rect 12440 38276 12492 38282
rect 12440 38218 12492 38224
rect 12452 37942 12480 38218
rect 12440 37936 12492 37942
rect 12440 37878 12492 37884
rect 12820 37874 12848 38286
rect 12256 37868 12308 37874
rect 12256 37810 12308 37816
rect 12808 37868 12860 37874
rect 12808 37810 12860 37816
rect 13556 37466 13584 39238
rect 13832 39098 13860 39306
rect 13912 39296 13964 39302
rect 13912 39238 13964 39244
rect 14004 39296 14056 39302
rect 14004 39238 14056 39244
rect 13924 39098 13952 39238
rect 13820 39092 13872 39098
rect 13820 39034 13872 39040
rect 13912 39092 13964 39098
rect 13912 39034 13964 39040
rect 13820 38752 13872 38758
rect 13820 38694 13872 38700
rect 13544 37460 13596 37466
rect 13544 37402 13596 37408
rect 13556 37330 13584 37402
rect 13544 37324 13596 37330
rect 13544 37266 13596 37272
rect 13832 37262 13860 38694
rect 13924 38332 13952 39034
rect 14016 39030 14044 39238
rect 14004 39024 14056 39030
rect 14004 38966 14056 38972
rect 14292 38486 14320 42350
rect 14464 40928 14516 40934
rect 14464 40870 14516 40876
rect 14476 40050 14504 40870
rect 14464 40044 14516 40050
rect 14464 39986 14516 39992
rect 14568 39574 14596 42706
rect 14648 42696 14700 42702
rect 14648 42638 14700 42644
rect 14660 41478 14688 42638
rect 14752 42226 14780 42842
rect 15016 42764 15068 42770
rect 15016 42706 15068 42712
rect 15028 42634 15056 42706
rect 15384 42696 15436 42702
rect 15384 42638 15436 42644
rect 15016 42628 15068 42634
rect 15016 42570 15068 42576
rect 15200 42356 15252 42362
rect 15200 42298 15252 42304
rect 14740 42220 14792 42226
rect 14740 42162 14792 42168
rect 15016 42084 15068 42090
rect 15016 42026 15068 42032
rect 15028 41818 15056 42026
rect 15016 41812 15068 41818
rect 15016 41754 15068 41760
rect 15212 41562 15240 42298
rect 15396 41750 15424 42638
rect 15580 41818 15608 43046
rect 15568 41812 15620 41818
rect 15568 41754 15620 41760
rect 15384 41744 15436 41750
rect 15384 41686 15436 41692
rect 15212 41534 15424 41562
rect 15396 41478 15424 41534
rect 14648 41472 14700 41478
rect 14648 41414 14700 41420
rect 15384 41472 15436 41478
rect 15384 41414 15436 41420
rect 14660 41206 14688 41414
rect 14648 41200 14700 41206
rect 14648 41142 14700 41148
rect 14556 39568 14608 39574
rect 14556 39510 14608 39516
rect 14280 38480 14332 38486
rect 14280 38422 14332 38428
rect 13924 38304 14044 38332
rect 14016 38214 14044 38304
rect 14004 38208 14056 38214
rect 14004 38150 14056 38156
rect 14292 37806 14320 38422
rect 14280 37800 14332 37806
rect 14280 37742 14332 37748
rect 14292 37398 14320 37742
rect 14280 37392 14332 37398
rect 14280 37334 14332 37340
rect 13820 37256 13872 37262
rect 13820 37198 13872 37204
rect 14568 36718 14596 39510
rect 14660 38282 14688 41142
rect 15200 40996 15252 41002
rect 15200 40938 15252 40944
rect 15292 40996 15344 41002
rect 15292 40938 15344 40944
rect 15212 40594 15240 40938
rect 15200 40588 15252 40594
rect 15200 40530 15252 40536
rect 15212 40050 15240 40530
rect 15200 40044 15252 40050
rect 15200 39986 15252 39992
rect 15108 39500 15160 39506
rect 15108 39442 15160 39448
rect 15120 38962 15148 39442
rect 15108 38956 15160 38962
rect 15108 38898 15160 38904
rect 14648 38276 14700 38282
rect 14648 38218 14700 38224
rect 14660 37942 14688 38218
rect 15120 38214 15148 38898
rect 15212 38554 15240 39986
rect 15304 39642 15332 40938
rect 15396 40526 15424 41414
rect 15672 41313 15700 43794
rect 16132 43314 16160 43930
rect 16396 43784 16448 43790
rect 16396 43726 16448 43732
rect 16120 43308 16172 43314
rect 16120 43250 16172 43256
rect 16028 43240 16080 43246
rect 16028 43182 16080 43188
rect 16040 42362 16068 43182
rect 16132 42770 16160 43250
rect 16212 43240 16264 43246
rect 16212 43182 16264 43188
rect 16224 42906 16252 43182
rect 16212 42900 16264 42906
rect 16212 42842 16264 42848
rect 16120 42764 16172 42770
rect 16120 42706 16172 42712
rect 16028 42356 16080 42362
rect 16028 42298 16080 42304
rect 16304 42084 16356 42090
rect 16304 42026 16356 42032
rect 15658 41304 15714 41313
rect 15658 41239 15660 41248
rect 15712 41239 15714 41248
rect 15660 41210 15712 41216
rect 16316 41002 16344 42026
rect 16408 41614 16436 43726
rect 16580 43172 16632 43178
rect 16580 43114 16632 43120
rect 16488 42356 16540 42362
rect 16488 42298 16540 42304
rect 16396 41608 16448 41614
rect 16396 41550 16448 41556
rect 16408 41478 16436 41550
rect 16396 41472 16448 41478
rect 16396 41414 16448 41420
rect 16304 40996 16356 41002
rect 16304 40938 16356 40944
rect 15384 40520 15436 40526
rect 15384 40462 15436 40468
rect 15292 39636 15344 39642
rect 15292 39578 15344 39584
rect 15396 39370 15424 40462
rect 15568 40384 15620 40390
rect 15568 40326 15620 40332
rect 15580 39642 15608 40326
rect 16316 39914 16344 40938
rect 16304 39908 16356 39914
rect 16304 39850 16356 39856
rect 16500 39642 16528 42298
rect 16592 41818 16620 43114
rect 16684 42838 16712 44390
rect 17328 43926 17356 44678
rect 21744 44538 21772 44746
rect 24032 44736 24084 44742
rect 24032 44678 24084 44684
rect 26606 44704 26662 44713
rect 20076 44532 20128 44538
rect 20076 44474 20128 44480
rect 21732 44532 21784 44538
rect 21732 44474 21784 44480
rect 17868 44396 17920 44402
rect 17868 44338 17920 44344
rect 17500 44192 17552 44198
rect 17500 44134 17552 44140
rect 17592 44192 17644 44198
rect 17592 44134 17644 44140
rect 17512 43926 17540 44134
rect 16856 43920 16908 43926
rect 16856 43862 16908 43868
rect 17316 43920 17368 43926
rect 17316 43862 17368 43868
rect 17500 43920 17552 43926
rect 17500 43862 17552 43868
rect 16868 43450 16896 43862
rect 16856 43444 16908 43450
rect 16856 43386 16908 43392
rect 16948 43444 17000 43450
rect 16948 43386 17000 43392
rect 16672 42832 16724 42838
rect 16672 42774 16724 42780
rect 16764 42696 16816 42702
rect 16764 42638 16816 42644
rect 16776 42362 16804 42638
rect 16764 42356 16816 42362
rect 16764 42298 16816 42304
rect 16868 42265 16896 43386
rect 16960 43178 16988 43386
rect 16948 43172 17000 43178
rect 16948 43114 17000 43120
rect 16960 42838 16988 43114
rect 16948 42832 17000 42838
rect 16948 42774 17000 42780
rect 16854 42256 16910 42265
rect 16672 42220 16724 42226
rect 16854 42191 16910 42200
rect 16672 42162 16724 42168
rect 16580 41812 16632 41818
rect 16580 41754 16632 41760
rect 16684 41682 16712 42162
rect 16960 42090 16988 42774
rect 17132 42560 17184 42566
rect 17132 42502 17184 42508
rect 17144 42158 17172 42502
rect 17132 42152 17184 42158
rect 17132 42094 17184 42100
rect 16948 42084 17000 42090
rect 16948 42026 17000 42032
rect 16672 41676 16724 41682
rect 16672 41618 16724 41624
rect 16764 41676 16816 41682
rect 16764 41618 16816 41624
rect 16776 41274 16804 41618
rect 16764 41268 16816 41274
rect 16764 41210 16816 41216
rect 16776 40662 16804 41210
rect 16948 40928 17000 40934
rect 16948 40870 17000 40876
rect 16960 40730 16988 40870
rect 16948 40724 17000 40730
rect 16948 40666 17000 40672
rect 16764 40656 16816 40662
rect 16764 40598 16816 40604
rect 16764 40520 16816 40526
rect 16764 40462 16816 40468
rect 15568 39636 15620 39642
rect 15568 39578 15620 39584
rect 16488 39636 16540 39642
rect 16488 39578 16540 39584
rect 16776 39438 16804 40462
rect 16856 40384 16908 40390
rect 16856 40326 16908 40332
rect 16868 40186 16896 40326
rect 16856 40180 16908 40186
rect 16856 40122 16908 40128
rect 17328 40050 17356 43862
rect 17512 43450 17540 43862
rect 17500 43444 17552 43450
rect 17500 43386 17552 43392
rect 17604 41818 17632 44134
rect 17880 42226 17908 44338
rect 18512 44328 18564 44334
rect 18512 44270 18564 44276
rect 19156 44328 19208 44334
rect 19208 44288 19288 44316
rect 19156 44270 19208 44276
rect 17958 43752 18014 43761
rect 17958 43687 17960 43696
rect 18012 43687 18014 43696
rect 17960 43658 18012 43664
rect 18052 43648 18104 43654
rect 18052 43590 18104 43596
rect 17960 42560 18012 42566
rect 17960 42502 18012 42508
rect 17868 42220 17920 42226
rect 17868 42162 17920 42168
rect 17684 42016 17736 42022
rect 17684 41958 17736 41964
rect 17696 41818 17724 41958
rect 17592 41812 17644 41818
rect 17592 41754 17644 41760
rect 17684 41812 17736 41818
rect 17684 41754 17736 41760
rect 17880 41614 17908 42162
rect 17972 42022 18000 42502
rect 18064 42226 18092 43590
rect 18524 43110 18552 44270
rect 18880 44260 18932 44266
rect 18880 44202 18932 44208
rect 18786 43480 18842 43489
rect 18786 43415 18842 43424
rect 18800 43382 18828 43415
rect 18788 43376 18840 43382
rect 18788 43318 18840 43324
rect 18892 43296 18920 44202
rect 18972 44192 19024 44198
rect 18972 44134 19024 44140
rect 18984 43926 19012 44134
rect 18972 43920 19024 43926
rect 18972 43862 19024 43868
rect 19260 43654 19288 44288
rect 19524 43852 19576 43858
rect 19524 43794 19576 43800
rect 19248 43648 19300 43654
rect 19248 43590 19300 43596
rect 19432 43648 19484 43654
rect 19432 43590 19484 43596
rect 19064 43308 19116 43314
rect 18892 43268 19064 43296
rect 19064 43250 19116 43256
rect 19260 43246 19288 43590
rect 19340 43308 19392 43314
rect 19340 43250 19392 43256
rect 19248 43240 19300 43246
rect 19248 43182 19300 43188
rect 18512 43104 18564 43110
rect 18512 43046 18564 43052
rect 19156 43104 19208 43110
rect 19156 43046 19208 43052
rect 19168 42226 19196 43046
rect 19352 42786 19380 43250
rect 19260 42758 19380 42786
rect 19260 42566 19288 42758
rect 19444 42702 19472 43590
rect 19536 42906 19564 43794
rect 19800 43784 19852 43790
rect 19798 43752 19800 43761
rect 19892 43784 19944 43790
rect 19852 43752 19854 43761
rect 19892 43726 19944 43732
rect 19798 43687 19854 43696
rect 19904 43450 19932 43726
rect 20088 43654 20116 44474
rect 20720 44260 20772 44266
rect 20720 44202 20772 44208
rect 20996 44260 21048 44266
rect 20996 44202 21048 44208
rect 21456 44260 21508 44266
rect 21456 44202 21508 44208
rect 20260 44192 20312 44198
rect 20260 44134 20312 44140
rect 20076 43648 20128 43654
rect 20076 43590 20128 43596
rect 19616 43444 19668 43450
rect 19616 43386 19668 43392
rect 19892 43444 19944 43450
rect 19892 43386 19944 43392
rect 19628 43314 19656 43386
rect 19616 43308 19668 43314
rect 19616 43250 19668 43256
rect 20088 43178 20116 43590
rect 20168 43308 20220 43314
rect 20168 43250 20220 43256
rect 20076 43172 20128 43178
rect 20076 43114 20128 43120
rect 20088 43058 20116 43114
rect 19904 43030 20116 43058
rect 19524 42900 19576 42906
rect 19524 42842 19576 42848
rect 19432 42696 19484 42702
rect 19432 42638 19484 42644
rect 19248 42560 19300 42566
rect 19248 42502 19300 42508
rect 19260 42226 19288 42502
rect 18052 42220 18104 42226
rect 18052 42162 18104 42168
rect 18420 42220 18472 42226
rect 18420 42162 18472 42168
rect 19156 42220 19208 42226
rect 19156 42162 19208 42168
rect 19248 42220 19300 42226
rect 19248 42162 19300 42168
rect 17960 42016 18012 42022
rect 17960 41958 18012 41964
rect 17972 41750 18000 41958
rect 17960 41744 18012 41750
rect 17960 41686 18012 41692
rect 17868 41608 17920 41614
rect 17868 41550 17920 41556
rect 18328 41608 18380 41614
rect 18328 41550 18380 41556
rect 17880 41138 17908 41550
rect 18052 41472 18104 41478
rect 18052 41414 18104 41420
rect 17500 41132 17552 41138
rect 17500 41074 17552 41080
rect 17868 41132 17920 41138
rect 17868 41074 17920 41080
rect 17960 41132 18012 41138
rect 17960 41074 18012 41080
rect 17408 40928 17460 40934
rect 17408 40870 17460 40876
rect 17420 40662 17448 40870
rect 17408 40656 17460 40662
rect 17408 40598 17460 40604
rect 17512 40526 17540 41074
rect 17972 40594 18000 41074
rect 18064 41070 18092 41414
rect 18052 41064 18104 41070
rect 18052 41006 18104 41012
rect 17960 40588 18012 40594
rect 17960 40530 18012 40536
rect 17500 40520 17552 40526
rect 17500 40462 17552 40468
rect 17776 40384 17828 40390
rect 17776 40326 17828 40332
rect 17316 40044 17368 40050
rect 17316 39986 17368 39992
rect 17328 39438 17356 39986
rect 17788 39574 17816 40326
rect 17972 40050 18000 40530
rect 18340 40526 18368 41550
rect 18432 40526 18460 42162
rect 18880 41540 18932 41546
rect 18880 41482 18932 41488
rect 18788 40996 18840 41002
rect 18788 40938 18840 40944
rect 18052 40520 18104 40526
rect 18052 40462 18104 40468
rect 18328 40520 18380 40526
rect 18328 40462 18380 40468
rect 18420 40520 18472 40526
rect 18420 40462 18472 40468
rect 17960 40044 18012 40050
rect 17960 39986 18012 39992
rect 17972 39642 18000 39986
rect 18064 39846 18092 40462
rect 18340 39914 18368 40462
rect 18328 39908 18380 39914
rect 18328 39850 18380 39856
rect 18052 39840 18104 39846
rect 18052 39782 18104 39788
rect 17960 39636 18012 39642
rect 17960 39578 18012 39584
rect 17776 39568 17828 39574
rect 17776 39510 17828 39516
rect 17500 39500 17552 39506
rect 17500 39442 17552 39448
rect 18052 39500 18104 39506
rect 18052 39442 18104 39448
rect 16764 39432 16816 39438
rect 16764 39374 16816 39380
rect 17316 39432 17368 39438
rect 17316 39374 17368 39380
rect 15384 39364 15436 39370
rect 15384 39306 15436 39312
rect 15396 38962 15424 39306
rect 16856 39296 16908 39302
rect 16856 39238 16908 39244
rect 15384 38956 15436 38962
rect 15384 38898 15436 38904
rect 15568 38888 15620 38894
rect 15568 38830 15620 38836
rect 15384 38752 15436 38758
rect 15384 38694 15436 38700
rect 15200 38548 15252 38554
rect 15200 38490 15252 38496
rect 15108 38208 15160 38214
rect 15108 38150 15160 38156
rect 14648 37936 14700 37942
rect 14648 37878 14700 37884
rect 15120 37874 15148 38150
rect 15212 37874 15240 38490
rect 15292 38344 15344 38350
rect 15292 38286 15344 38292
rect 15108 37868 15160 37874
rect 15108 37810 15160 37816
rect 15200 37868 15252 37874
rect 15200 37810 15252 37816
rect 14830 37768 14886 37777
rect 14830 37703 14886 37712
rect 14556 36712 14608 36718
rect 14556 36654 14608 36660
rect 12162 36000 12218 36009
rect 12162 35935 12218 35944
rect 14844 35766 14872 37703
rect 15016 37664 15068 37670
rect 15016 37606 15068 37612
rect 8208 35760 8260 35766
rect 8206 35728 8208 35737
rect 14832 35760 14884 35766
rect 8260 35728 8262 35737
rect 15028 35737 15056 37606
rect 15120 37482 15148 37810
rect 15120 37454 15240 37482
rect 15106 37360 15162 37369
rect 15106 37295 15162 37304
rect 15120 36689 15148 37295
rect 15106 36680 15162 36689
rect 15212 36666 15240 37454
rect 15304 37262 15332 38286
rect 15396 38010 15424 38694
rect 15580 38554 15608 38830
rect 16212 38820 16264 38826
rect 16212 38762 16264 38768
rect 15568 38548 15620 38554
rect 15568 38490 15620 38496
rect 16224 38486 16252 38762
rect 16396 38752 16448 38758
rect 16396 38694 16448 38700
rect 16212 38480 16264 38486
rect 16212 38422 16264 38428
rect 16120 38208 16172 38214
rect 16120 38150 16172 38156
rect 16132 38010 16160 38150
rect 15384 38004 15436 38010
rect 15384 37946 15436 37952
rect 16120 38004 16172 38010
rect 16120 37946 16172 37952
rect 16224 37806 16252 38422
rect 16408 38350 16436 38694
rect 16396 38344 16448 38350
rect 16396 38286 16448 38292
rect 16212 37800 16264 37806
rect 16212 37742 16264 37748
rect 16868 37262 16896 39238
rect 17512 39098 17540 39442
rect 17500 39092 17552 39098
rect 17500 39034 17552 39040
rect 17224 38412 17276 38418
rect 17224 38354 17276 38360
rect 17236 38010 17264 38354
rect 17684 38344 17736 38350
rect 17684 38286 17736 38292
rect 17224 38004 17276 38010
rect 17224 37946 17276 37952
rect 17236 37466 17264 37946
rect 17696 37466 17724 38286
rect 18064 37942 18092 39442
rect 18432 39370 18460 40462
rect 18512 39840 18564 39846
rect 18512 39782 18564 39788
rect 18420 39364 18472 39370
rect 18420 39306 18472 39312
rect 18524 39030 18552 39782
rect 18800 39574 18828 40938
rect 18788 39568 18840 39574
rect 18788 39510 18840 39516
rect 18512 39024 18564 39030
rect 18512 38966 18564 38972
rect 18800 38570 18828 39510
rect 18892 39438 18920 41482
rect 19616 41472 19668 41478
rect 19154 41440 19210 41449
rect 19616 41414 19668 41420
rect 19904 41414 19932 43030
rect 19984 42900 20036 42906
rect 19984 42842 20036 42848
rect 19154 41375 19210 41384
rect 19168 41206 19196 41375
rect 19156 41200 19208 41206
rect 19156 41142 19208 41148
rect 19064 41064 19116 41070
rect 19064 41006 19116 41012
rect 19076 39846 19104 41006
rect 19340 40520 19392 40526
rect 19340 40462 19392 40468
rect 19064 39840 19116 39846
rect 19064 39782 19116 39788
rect 19156 39840 19208 39846
rect 19156 39782 19208 39788
rect 19076 39574 19104 39782
rect 19168 39642 19196 39782
rect 19156 39636 19208 39642
rect 19156 39578 19208 39584
rect 19064 39568 19116 39574
rect 19064 39510 19116 39516
rect 18880 39432 18932 39438
rect 18880 39374 18932 39380
rect 18708 38542 18828 38570
rect 18144 38480 18196 38486
rect 18144 38422 18196 38428
rect 18052 37936 18104 37942
rect 18052 37878 18104 37884
rect 17224 37460 17276 37466
rect 17224 37402 17276 37408
rect 17684 37460 17736 37466
rect 17684 37402 17736 37408
rect 18156 37398 18184 38422
rect 18708 37806 18736 38542
rect 18696 37800 18748 37806
rect 18696 37742 18748 37748
rect 18144 37392 18196 37398
rect 18144 37334 18196 37340
rect 18892 37262 18920 39374
rect 19352 39098 19380 40462
rect 19340 39092 19392 39098
rect 19340 39034 19392 39040
rect 19628 38894 19656 41414
rect 19812 41386 19932 41414
rect 19812 40186 19840 41386
rect 19996 41138 20024 42842
rect 20180 42838 20208 43250
rect 20272 42906 20300 44134
rect 20732 44010 20760 44202
rect 20640 43982 20760 44010
rect 20640 43790 20668 43982
rect 20720 43920 20772 43926
rect 20720 43862 20772 43868
rect 20628 43784 20680 43790
rect 20628 43726 20680 43732
rect 20732 43314 20760 43862
rect 20812 43852 20864 43858
rect 20812 43794 20864 43800
rect 20720 43308 20772 43314
rect 20720 43250 20772 43256
rect 20260 42900 20312 42906
rect 20260 42842 20312 42848
rect 20168 42832 20220 42838
rect 20168 42774 20220 42780
rect 19984 41132 20036 41138
rect 19984 41074 20036 41080
rect 19892 40520 19944 40526
rect 19892 40462 19944 40468
rect 19800 40180 19852 40186
rect 19800 40122 19852 40128
rect 19904 39914 19932 40462
rect 19996 40066 20024 41074
rect 20180 41018 20208 42774
rect 20732 42362 20760 43250
rect 20824 42906 20852 43794
rect 20812 42900 20864 42906
rect 20812 42842 20864 42848
rect 20904 42764 20956 42770
rect 20904 42706 20956 42712
rect 20812 42560 20864 42566
rect 20812 42502 20864 42508
rect 20824 42362 20852 42502
rect 20720 42356 20772 42362
rect 20720 42298 20772 42304
rect 20812 42356 20864 42362
rect 20812 42298 20864 42304
rect 20536 42084 20588 42090
rect 20536 42026 20588 42032
rect 20260 41472 20312 41478
rect 20260 41414 20312 41420
rect 20272 41138 20300 41414
rect 20260 41132 20312 41138
rect 20260 41074 20312 41080
rect 20180 41002 20392 41018
rect 20180 40996 20404 41002
rect 20180 40990 20352 40996
rect 20352 40938 20404 40944
rect 20364 40526 20392 40938
rect 20444 40588 20496 40594
rect 20444 40530 20496 40536
rect 20352 40520 20404 40526
rect 20352 40462 20404 40468
rect 20456 40186 20484 40530
rect 20444 40180 20496 40186
rect 20444 40122 20496 40128
rect 19996 40050 20116 40066
rect 19996 40044 20128 40050
rect 19996 40038 20076 40044
rect 20076 39986 20128 39992
rect 19892 39908 19944 39914
rect 19892 39850 19944 39856
rect 20088 39642 20116 39986
rect 20076 39636 20128 39642
rect 20076 39578 20128 39584
rect 19984 39364 20036 39370
rect 19984 39306 20036 39312
rect 19892 39296 19944 39302
rect 19892 39238 19944 39244
rect 19708 39092 19760 39098
rect 19708 39034 19760 39040
rect 19432 38888 19484 38894
rect 19432 38830 19484 38836
rect 19616 38888 19668 38894
rect 19616 38830 19668 38836
rect 19340 38344 19392 38350
rect 19340 38286 19392 38292
rect 19064 38208 19116 38214
rect 19248 38208 19300 38214
rect 19116 38156 19196 38162
rect 19064 38150 19196 38156
rect 19248 38150 19300 38156
rect 19076 38134 19196 38150
rect 19168 37806 19196 38134
rect 19156 37800 19208 37806
rect 19156 37742 19208 37748
rect 15292 37256 15344 37262
rect 15292 37198 15344 37204
rect 16856 37256 16908 37262
rect 16856 37198 16908 37204
rect 18880 37256 18932 37262
rect 18880 37198 18932 37204
rect 19168 36786 19196 37742
rect 19260 37738 19288 38150
rect 19352 38010 19380 38286
rect 19340 38004 19392 38010
rect 19340 37946 19392 37952
rect 19248 37732 19300 37738
rect 19248 37674 19300 37680
rect 19260 37398 19288 37674
rect 19444 37466 19472 38830
rect 19522 38720 19578 38729
rect 19522 38655 19578 38664
rect 19432 37460 19484 37466
rect 19432 37402 19484 37408
rect 19248 37392 19300 37398
rect 19248 37334 19300 37340
rect 19536 37097 19564 38655
rect 19522 37088 19578 37097
rect 19522 37023 19578 37032
rect 19156 36780 19208 36786
rect 19156 36722 19208 36728
rect 15290 36680 15346 36689
rect 15212 36638 15290 36666
rect 15106 36615 15162 36624
rect 15290 36615 15346 36624
rect 19720 36009 19748 39034
rect 19904 38962 19932 39238
rect 19996 38962 20024 39306
rect 19892 38956 19944 38962
rect 19892 38898 19944 38904
rect 19984 38956 20036 38962
rect 19984 38898 20036 38904
rect 20260 38752 20312 38758
rect 20260 38694 20312 38700
rect 20352 38752 20404 38758
rect 20352 38694 20404 38700
rect 20272 38350 20300 38694
rect 20260 38344 20312 38350
rect 20260 38286 20312 38292
rect 20364 36961 20392 38694
rect 20456 38554 20484 40122
rect 20548 38826 20576 42026
rect 20732 41818 20760 42298
rect 20720 41812 20772 41818
rect 20720 41754 20772 41760
rect 20628 41608 20680 41614
rect 20628 41550 20680 41556
rect 20640 40390 20668 41550
rect 20732 41414 20760 41754
rect 20732 41386 20852 41414
rect 20824 40730 20852 41386
rect 20916 40905 20944 42706
rect 21008 41614 21036 44202
rect 21468 42702 21496 44202
rect 21548 44192 21600 44198
rect 21548 44134 21600 44140
rect 21560 43926 21588 44134
rect 21548 43920 21600 43926
rect 21548 43862 21600 43868
rect 21744 43246 21772 44474
rect 22284 44396 22336 44402
rect 22284 44338 22336 44344
rect 23940 44396 23992 44402
rect 23940 44338 23992 44344
rect 22100 44192 22152 44198
rect 22100 44134 22152 44140
rect 21916 43648 21968 43654
rect 21916 43590 21968 43596
rect 21928 43450 21956 43590
rect 22112 43450 22140 44134
rect 22192 43920 22244 43926
rect 22192 43862 22244 43868
rect 21916 43444 21968 43450
rect 21916 43386 21968 43392
rect 22100 43444 22152 43450
rect 22100 43386 22152 43392
rect 21732 43240 21784 43246
rect 21732 43182 21784 43188
rect 21928 43092 21956 43386
rect 22100 43172 22152 43178
rect 22100 43114 22152 43120
rect 22008 43104 22060 43110
rect 21928 43064 22008 43092
rect 22008 43046 22060 43052
rect 22112 42838 22140 43114
rect 22204 43110 22232 43862
rect 22296 43790 22324 44338
rect 22560 44328 22612 44334
rect 22560 44270 22612 44276
rect 22468 44192 22520 44198
rect 22468 44134 22520 44140
rect 22284 43784 22336 43790
rect 22284 43726 22336 43732
rect 22480 43314 22508 44134
rect 22468 43308 22520 43314
rect 22468 43250 22520 43256
rect 22192 43104 22244 43110
rect 22192 43046 22244 43052
rect 22100 42832 22152 42838
rect 22100 42774 22152 42780
rect 21456 42696 21508 42702
rect 21456 42638 21508 42644
rect 20996 41608 21048 41614
rect 20996 41550 21048 41556
rect 21008 41414 21036 41550
rect 21272 41540 21324 41546
rect 21272 41482 21324 41488
rect 21008 41386 21128 41414
rect 20996 41268 21048 41274
rect 20996 41210 21048 41216
rect 20902 40896 20958 40905
rect 20902 40831 20958 40840
rect 20812 40724 20864 40730
rect 20812 40666 20864 40672
rect 20720 40520 20772 40526
rect 20720 40462 20772 40468
rect 20628 40384 20680 40390
rect 20628 40326 20680 40332
rect 20640 39506 20668 40326
rect 20628 39500 20680 39506
rect 20628 39442 20680 39448
rect 20732 39386 20760 40462
rect 21008 39982 21036 41210
rect 21100 40118 21128 41386
rect 21284 40730 21312 41482
rect 21468 41138 21496 42638
rect 22100 42356 22152 42362
rect 22100 42298 22152 42304
rect 21824 42220 21876 42226
rect 21824 42162 21876 42168
rect 21548 41608 21600 41614
rect 21548 41550 21600 41556
rect 21560 41274 21588 41550
rect 21732 41472 21784 41478
rect 21732 41414 21784 41420
rect 21548 41268 21600 41274
rect 21548 41210 21600 41216
rect 21744 41206 21772 41414
rect 21732 41200 21784 41206
rect 21732 41142 21784 41148
rect 21456 41132 21508 41138
rect 21456 41074 21508 41080
rect 21272 40724 21324 40730
rect 21272 40666 21324 40672
rect 21468 40526 21496 41074
rect 21456 40520 21508 40526
rect 21456 40462 21508 40468
rect 21640 40452 21692 40458
rect 21640 40394 21692 40400
rect 21652 40118 21680 40394
rect 21088 40112 21140 40118
rect 21088 40054 21140 40060
rect 21640 40112 21692 40118
rect 21640 40054 21692 40060
rect 20996 39976 21048 39982
rect 20996 39918 21048 39924
rect 21548 39636 21600 39642
rect 21548 39578 21600 39584
rect 20640 39370 20760 39386
rect 21364 39432 21416 39438
rect 21364 39374 21416 39380
rect 20628 39364 20760 39370
rect 20680 39358 20760 39364
rect 20812 39364 20864 39370
rect 20628 39306 20680 39312
rect 20812 39306 20864 39312
rect 20628 38956 20680 38962
rect 20628 38898 20680 38904
rect 20536 38820 20588 38826
rect 20536 38762 20588 38768
rect 20444 38548 20496 38554
rect 20444 38490 20496 38496
rect 20640 37466 20668 38898
rect 20824 38842 20852 39306
rect 21376 38962 21404 39374
rect 21364 38956 21416 38962
rect 21364 38898 21416 38904
rect 20732 38814 20852 38842
rect 21088 38888 21140 38894
rect 21088 38830 21140 38836
rect 20732 38758 20760 38814
rect 20720 38752 20772 38758
rect 20720 38694 20772 38700
rect 20812 38752 20864 38758
rect 20812 38694 20864 38700
rect 20824 37738 20852 38694
rect 21100 38554 21128 38830
rect 20904 38548 20956 38554
rect 20904 38490 20956 38496
rect 21088 38548 21140 38554
rect 21088 38490 21140 38496
rect 20916 37738 20944 38490
rect 21560 38418 21588 39578
rect 21640 39500 21692 39506
rect 21640 39442 21692 39448
rect 21548 38412 21600 38418
rect 21548 38354 21600 38360
rect 20720 37732 20772 37738
rect 20720 37674 20772 37680
rect 20812 37732 20864 37738
rect 20812 37674 20864 37680
rect 20904 37732 20956 37738
rect 20904 37674 20956 37680
rect 20628 37460 20680 37466
rect 20628 37402 20680 37408
rect 20732 37262 20760 37674
rect 20720 37256 20772 37262
rect 21652 37233 21680 39442
rect 21836 39438 21864 42162
rect 22112 40508 22140 42298
rect 22204 41750 22232 43046
rect 22572 42906 22600 44270
rect 23388 44260 23440 44266
rect 23388 44202 23440 44208
rect 23400 43858 23428 44202
rect 22836 43852 22888 43858
rect 22836 43794 22888 43800
rect 23388 43852 23440 43858
rect 23388 43794 23440 43800
rect 22744 43784 22796 43790
rect 22744 43726 22796 43732
rect 22652 43648 22704 43654
rect 22652 43590 22704 43596
rect 22664 43314 22692 43590
rect 22652 43308 22704 43314
rect 22652 43250 22704 43256
rect 22560 42900 22612 42906
rect 22560 42842 22612 42848
rect 22376 42764 22428 42770
rect 22376 42706 22428 42712
rect 22388 42566 22416 42706
rect 22560 42696 22612 42702
rect 22560 42638 22612 42644
rect 22376 42560 22428 42566
rect 22376 42502 22428 42508
rect 22388 42022 22416 42502
rect 22572 42226 22600 42638
rect 22664 42362 22692 43250
rect 22756 42906 22784 43726
rect 22744 42900 22796 42906
rect 22744 42842 22796 42848
rect 22848 42702 22876 43794
rect 23952 43450 23980 44338
rect 24044 44334 24072 44678
rect 26606 44639 26662 44648
rect 26424 44464 26476 44470
rect 26238 44432 26294 44441
rect 26424 44406 26476 44412
rect 26238 44367 26294 44376
rect 26252 44334 26280 44367
rect 24032 44328 24084 44334
rect 24032 44270 24084 44276
rect 26240 44328 26292 44334
rect 26240 44270 26292 44276
rect 26056 44260 26108 44266
rect 26056 44202 26108 44208
rect 25044 44192 25096 44198
rect 25044 44134 25096 44140
rect 25320 44192 25372 44198
rect 25504 44192 25556 44198
rect 25320 44134 25372 44140
rect 25424 44152 25504 44180
rect 24124 43988 24176 43994
rect 24124 43930 24176 43936
rect 23940 43444 23992 43450
rect 23940 43386 23992 43392
rect 23572 43376 23624 43382
rect 23624 43324 23704 43330
rect 23572 43318 23704 43324
rect 23584 43302 23704 43318
rect 23676 43246 23704 43302
rect 24136 43246 24164 43930
rect 24952 43920 25004 43926
rect 24952 43862 25004 43868
rect 24584 43716 24636 43722
rect 24584 43658 24636 43664
rect 24596 43314 24624 43658
rect 24584 43308 24636 43314
rect 24584 43250 24636 43256
rect 23664 43240 23716 43246
rect 23664 43182 23716 43188
rect 24124 43240 24176 43246
rect 24124 43182 24176 43188
rect 24964 43178 24992 43862
rect 23848 43172 23900 43178
rect 23848 43114 23900 43120
rect 24584 43172 24636 43178
rect 24584 43114 24636 43120
rect 24952 43172 25004 43178
rect 24952 43114 25004 43120
rect 22928 43104 22980 43110
rect 22928 43046 22980 43052
rect 22836 42696 22888 42702
rect 22836 42638 22888 42644
rect 22652 42356 22704 42362
rect 22652 42298 22704 42304
rect 22560 42220 22612 42226
rect 22560 42162 22612 42168
rect 22940 42158 22968 43046
rect 23388 42696 23440 42702
rect 23388 42638 23440 42644
rect 23112 42288 23164 42294
rect 23112 42230 23164 42236
rect 23204 42288 23256 42294
rect 23204 42230 23256 42236
rect 23020 42220 23072 42226
rect 23020 42162 23072 42168
rect 22928 42152 22980 42158
rect 22928 42094 22980 42100
rect 22376 42016 22428 42022
rect 22376 41958 22428 41964
rect 22192 41744 22244 41750
rect 22192 41686 22244 41692
rect 22388 41585 22416 41958
rect 22836 41608 22888 41614
rect 22374 41576 22430 41585
rect 22836 41550 22888 41556
rect 22374 41511 22430 41520
rect 22560 41200 22612 41206
rect 22560 41142 22612 41148
rect 22192 40928 22244 40934
rect 22192 40870 22244 40876
rect 22284 40928 22336 40934
rect 22284 40870 22336 40876
rect 22204 40730 22232 40870
rect 22192 40724 22244 40730
rect 22192 40666 22244 40672
rect 22192 40520 22244 40526
rect 22112 40480 22192 40508
rect 22192 40462 22244 40468
rect 22100 40384 22152 40390
rect 22100 40326 22152 40332
rect 22112 40050 22140 40326
rect 22204 40118 22232 40462
rect 22296 40186 22324 40870
rect 22284 40180 22336 40186
rect 22284 40122 22336 40128
rect 22192 40112 22244 40118
rect 22192 40054 22244 40060
rect 22572 40050 22600 41142
rect 22848 40594 22876 41550
rect 23032 41070 23060 42162
rect 23124 41478 23152 42230
rect 23216 42022 23244 42230
rect 23204 42016 23256 42022
rect 23204 41958 23256 41964
rect 23400 41750 23428 42638
rect 23480 42560 23532 42566
rect 23480 42502 23532 42508
rect 23492 41818 23520 42502
rect 23860 41818 23888 43114
rect 24216 42900 24268 42906
rect 24216 42842 24268 42848
rect 24228 42158 24256 42842
rect 24596 42362 24624 43114
rect 24964 42838 24992 43114
rect 24952 42832 25004 42838
rect 24952 42774 25004 42780
rect 24676 42628 24728 42634
rect 24676 42570 24728 42576
rect 24584 42356 24636 42362
rect 24584 42298 24636 42304
rect 24216 42152 24268 42158
rect 24216 42094 24268 42100
rect 24584 42152 24636 42158
rect 24584 42094 24636 42100
rect 24124 42016 24176 42022
rect 24124 41958 24176 41964
rect 24216 42016 24268 42022
rect 24216 41958 24268 41964
rect 23480 41812 23532 41818
rect 23480 41754 23532 41760
rect 23664 41812 23716 41818
rect 23664 41754 23716 41760
rect 23848 41812 23900 41818
rect 23848 41754 23900 41760
rect 23388 41744 23440 41750
rect 23388 41686 23440 41692
rect 23112 41472 23164 41478
rect 23112 41414 23164 41420
rect 23020 41064 23072 41070
rect 23020 41006 23072 41012
rect 22836 40588 22888 40594
rect 22836 40530 22888 40536
rect 23676 40526 23704 41754
rect 23860 41682 23888 41754
rect 24030 41712 24086 41721
rect 23848 41676 23900 41682
rect 24030 41647 24086 41656
rect 23848 41618 23900 41624
rect 23756 41608 23808 41614
rect 23756 41550 23808 41556
rect 23768 41274 23796 41550
rect 23756 41268 23808 41274
rect 23756 41210 23808 41216
rect 23940 40656 23992 40662
rect 23940 40598 23992 40604
rect 23572 40520 23624 40526
rect 23572 40462 23624 40468
rect 23664 40520 23716 40526
rect 23664 40462 23716 40468
rect 22928 40384 22980 40390
rect 22928 40326 22980 40332
rect 23296 40384 23348 40390
rect 23296 40326 23348 40332
rect 22100 40044 22152 40050
rect 22100 39986 22152 39992
rect 22560 40044 22612 40050
rect 22560 39986 22612 39992
rect 22940 39982 22968 40326
rect 23308 40118 23336 40326
rect 23296 40112 23348 40118
rect 23296 40054 23348 40060
rect 22928 39976 22980 39982
rect 22928 39918 22980 39924
rect 22744 39840 22796 39846
rect 22744 39782 22796 39788
rect 22756 39574 22784 39782
rect 22744 39568 22796 39574
rect 22744 39510 22796 39516
rect 21824 39432 21876 39438
rect 21824 39374 21876 39380
rect 21836 38842 21864 39374
rect 21836 38814 21956 38842
rect 21824 38752 21876 38758
rect 21824 38694 21876 38700
rect 21836 37466 21864 38694
rect 21824 37460 21876 37466
rect 21824 37402 21876 37408
rect 21836 37330 21864 37402
rect 21824 37324 21876 37330
rect 21824 37266 21876 37272
rect 21928 37262 21956 38814
rect 23204 38820 23256 38826
rect 23204 38762 23256 38768
rect 23020 38752 23072 38758
rect 23020 38694 23072 38700
rect 22836 38344 22888 38350
rect 22836 38286 22888 38292
rect 22848 37942 22876 38286
rect 22836 37936 22888 37942
rect 22836 37878 22888 37884
rect 23032 37806 23060 38694
rect 23020 37800 23072 37806
rect 23020 37742 23072 37748
rect 22284 37664 22336 37670
rect 22284 37606 22336 37612
rect 22296 37330 22324 37606
rect 22284 37324 22336 37330
rect 22284 37266 22336 37272
rect 21916 37256 21968 37262
rect 20720 37198 20772 37204
rect 21638 37224 21694 37233
rect 21916 37198 21968 37204
rect 21638 37159 21694 37168
rect 20350 36952 20406 36961
rect 20350 36887 20406 36896
rect 21638 36952 21694 36961
rect 21638 36887 21694 36896
rect 21652 36378 21680 36887
rect 23216 36825 23244 38762
rect 23308 37942 23336 40054
rect 23584 39982 23612 40462
rect 23572 39976 23624 39982
rect 23572 39918 23624 39924
rect 23480 38888 23532 38894
rect 23480 38830 23532 38836
rect 23492 38554 23520 38830
rect 23480 38548 23532 38554
rect 23480 38490 23532 38496
rect 23676 38350 23704 40462
rect 23952 40186 23980 40598
rect 23940 40180 23992 40186
rect 23940 40122 23992 40128
rect 23756 38752 23808 38758
rect 23756 38694 23808 38700
rect 23768 38486 23796 38694
rect 23756 38480 23808 38486
rect 23756 38422 23808 38428
rect 23664 38344 23716 38350
rect 23664 38286 23716 38292
rect 23480 38208 23532 38214
rect 23480 38150 23532 38156
rect 23296 37936 23348 37942
rect 23296 37878 23348 37884
rect 23388 37868 23440 37874
rect 23492 37856 23520 38150
rect 23440 37828 23520 37856
rect 23388 37810 23440 37816
rect 23848 37664 23900 37670
rect 23848 37606 23900 37612
rect 23860 37466 23888 37606
rect 23848 37460 23900 37466
rect 23848 37402 23900 37408
rect 23202 36816 23258 36825
rect 23202 36751 23258 36760
rect 22008 36644 22060 36650
rect 22008 36586 22060 36592
rect 21640 36372 21692 36378
rect 21640 36314 21692 36320
rect 19706 36000 19762 36009
rect 19706 35935 19762 35944
rect 20076 35964 20128 35970
rect 20076 35906 20128 35912
rect 20088 35737 20116 35906
rect 21364 35896 21416 35902
rect 22020 35873 22048 36586
rect 23204 36304 23256 36310
rect 24044 36281 24072 41647
rect 24136 41614 24164 41958
rect 24228 41750 24256 41958
rect 24216 41744 24268 41750
rect 24216 41686 24268 41692
rect 24124 41608 24176 41614
rect 24124 41550 24176 41556
rect 24596 41018 24624 42094
rect 24688 41138 24716 42570
rect 24964 42514 24992 42774
rect 24872 42486 24992 42514
rect 24768 42288 24820 42294
rect 24768 42230 24820 42236
rect 24676 41132 24728 41138
rect 24676 41074 24728 41080
rect 24780 41070 24808 42230
rect 24872 41750 24900 42486
rect 25056 42226 25084 44134
rect 25332 43790 25360 44134
rect 25320 43784 25372 43790
rect 25320 43726 25372 43732
rect 25332 43110 25360 43726
rect 25136 43104 25188 43110
rect 25136 43046 25188 43052
rect 25320 43104 25372 43110
rect 25320 43046 25372 43052
rect 25148 42362 25176 43046
rect 25424 42906 25452 44152
rect 25504 44134 25556 44140
rect 25596 44192 25648 44198
rect 25596 44134 25648 44140
rect 25608 43450 25636 44134
rect 25964 43784 26016 43790
rect 25964 43726 26016 43732
rect 25976 43450 26004 43726
rect 25596 43444 25648 43450
rect 25596 43386 25648 43392
rect 25964 43444 26016 43450
rect 25964 43386 26016 43392
rect 25504 43376 25556 43382
rect 25504 43318 25556 43324
rect 25412 42900 25464 42906
rect 25412 42842 25464 42848
rect 25136 42356 25188 42362
rect 25136 42298 25188 42304
rect 25044 42220 25096 42226
rect 25044 42162 25096 42168
rect 24860 41744 24912 41750
rect 24860 41686 24912 41692
rect 24872 41414 24900 41686
rect 25148 41614 25176 42298
rect 25412 42016 25464 42022
rect 25516 41970 25544 43318
rect 25872 42764 25924 42770
rect 25872 42706 25924 42712
rect 25780 42084 25832 42090
rect 25780 42026 25832 42032
rect 25464 41964 25544 41970
rect 25412 41958 25544 41964
rect 25424 41942 25544 41958
rect 25792 41818 25820 42026
rect 25884 42022 25912 42706
rect 26068 42702 26096 44202
rect 26240 43988 26292 43994
rect 26240 43930 26292 43936
rect 26252 43858 26280 43930
rect 26240 43852 26292 43858
rect 26240 43794 26292 43800
rect 26332 43784 26384 43790
rect 26160 43732 26332 43738
rect 26160 43726 26384 43732
rect 26160 43710 26372 43726
rect 26160 43110 26188 43710
rect 26240 43648 26292 43654
rect 26240 43590 26292 43596
rect 26252 43382 26280 43590
rect 26240 43376 26292 43382
rect 26240 43318 26292 43324
rect 26332 43376 26384 43382
rect 26332 43318 26384 43324
rect 26148 43104 26200 43110
rect 26148 43046 26200 43052
rect 26160 42906 26188 43046
rect 26148 42900 26200 42906
rect 26148 42842 26200 42848
rect 26056 42696 26108 42702
rect 26056 42638 26108 42644
rect 25964 42220 26016 42226
rect 26068 42208 26096 42638
rect 26240 42220 26292 42226
rect 26068 42180 26240 42208
rect 25964 42162 26016 42168
rect 26240 42162 26292 42168
rect 25976 42106 26004 42162
rect 26344 42106 26372 43318
rect 26436 42770 26464 44406
rect 26620 44334 26648 44639
rect 26790 44432 26846 44441
rect 26790 44367 26792 44376
rect 26844 44367 26846 44376
rect 27526 44432 27582 44441
rect 27526 44367 27528 44376
rect 26792 44338 26844 44344
rect 27580 44367 27582 44376
rect 27528 44338 27580 44344
rect 26608 44328 26660 44334
rect 26608 44270 26660 44276
rect 27436 44328 27488 44334
rect 27436 44270 27488 44276
rect 27344 44192 27396 44198
rect 27344 44134 27396 44140
rect 26884 43988 26936 43994
rect 26884 43930 26936 43936
rect 26514 43752 26570 43761
rect 26514 43687 26570 43696
rect 26528 43654 26556 43687
rect 26516 43648 26568 43654
rect 26516 43590 26568 43596
rect 26516 43104 26568 43110
rect 26516 43046 26568 43052
rect 26528 42906 26556 43046
rect 26516 42900 26568 42906
rect 26516 42842 26568 42848
rect 26424 42764 26476 42770
rect 26424 42706 26476 42712
rect 26606 42664 26662 42673
rect 26606 42599 26608 42608
rect 26660 42599 26662 42608
rect 26608 42570 26660 42576
rect 26700 42560 26752 42566
rect 26700 42502 26752 42508
rect 25976 42078 26372 42106
rect 25872 42016 25924 42022
rect 25872 41958 25924 41964
rect 25780 41812 25832 41818
rect 25780 41754 25832 41760
rect 26240 41676 26292 41682
rect 26240 41618 26292 41624
rect 25136 41608 25188 41614
rect 25136 41550 25188 41556
rect 25872 41540 25924 41546
rect 25872 41482 25924 41488
rect 24872 41386 25268 41414
rect 25240 41206 25268 41386
rect 25596 41268 25648 41274
rect 25596 41210 25648 41216
rect 25228 41200 25280 41206
rect 25228 41142 25280 41148
rect 25136 41132 25188 41138
rect 25136 41074 25188 41080
rect 24768 41064 24820 41070
rect 24596 40990 24716 41018
rect 24768 41006 24820 41012
rect 24688 40934 24716 40990
rect 24400 40928 24452 40934
rect 24400 40870 24452 40876
rect 24676 40928 24728 40934
rect 24676 40870 24728 40876
rect 24860 40928 24912 40934
rect 24860 40870 24912 40876
rect 24412 40050 24440 40870
rect 24768 40724 24820 40730
rect 24768 40666 24820 40672
rect 24492 40112 24544 40118
rect 24492 40054 24544 40060
rect 24400 40044 24452 40050
rect 24400 39986 24452 39992
rect 24216 39976 24268 39982
rect 24216 39918 24268 39924
rect 24228 39438 24256 39918
rect 24216 39432 24268 39438
rect 24216 39374 24268 39380
rect 24124 39024 24176 39030
rect 24124 38966 24176 38972
rect 24136 38729 24164 38966
rect 24504 38962 24532 40054
rect 24676 39840 24728 39846
rect 24676 39782 24728 39788
rect 24688 39030 24716 39782
rect 24780 39574 24808 40666
rect 24872 40633 24900 40870
rect 24858 40624 24914 40633
rect 24858 40559 24914 40568
rect 25148 40526 25176 41074
rect 25240 40662 25268 41142
rect 25502 41032 25558 41041
rect 25502 40967 25558 40976
rect 25228 40656 25280 40662
rect 25228 40598 25280 40604
rect 25136 40520 25188 40526
rect 25136 40462 25188 40468
rect 24952 39908 25004 39914
rect 24952 39850 25004 39856
rect 24768 39568 24820 39574
rect 24768 39510 24820 39516
rect 24964 39030 24992 39850
rect 25044 39636 25096 39642
rect 25044 39578 25096 39584
rect 24676 39024 24728 39030
rect 24676 38966 24728 38972
rect 24952 39024 25004 39030
rect 24952 38966 25004 38972
rect 24492 38956 24544 38962
rect 24492 38898 24544 38904
rect 25056 38894 25084 39578
rect 25240 39438 25268 40598
rect 25412 39976 25464 39982
rect 25412 39918 25464 39924
rect 25228 39432 25280 39438
rect 25228 39374 25280 39380
rect 25136 38956 25188 38962
rect 25136 38898 25188 38904
rect 25044 38888 25096 38894
rect 25044 38830 25096 38836
rect 24122 38720 24178 38729
rect 24122 38655 24178 38664
rect 25148 38593 25176 38898
rect 25134 38584 25190 38593
rect 25134 38519 25136 38528
rect 25188 38519 25190 38528
rect 25136 38490 25188 38496
rect 25148 37466 25176 38490
rect 25424 38418 25452 39918
rect 25412 38412 25464 38418
rect 25412 38354 25464 38360
rect 25424 37738 25452 38354
rect 25412 37732 25464 37738
rect 25412 37674 25464 37680
rect 25136 37460 25188 37466
rect 25136 37402 25188 37408
rect 24308 37324 24360 37330
rect 24308 37266 24360 37272
rect 23204 36246 23256 36252
rect 24030 36272 24086 36281
rect 21364 35838 21416 35844
rect 22006 35864 22062 35873
rect 21376 35737 21404 35838
rect 22006 35799 22062 35808
rect 23216 35737 23244 36246
rect 24030 36207 24086 36216
rect 23572 36168 23624 36174
rect 23572 36110 23624 36116
rect 23584 35873 23612 36110
rect 24320 35970 24348 37266
rect 24768 36916 24820 36922
rect 24768 36858 24820 36864
rect 24780 36825 24808 36858
rect 24766 36816 24822 36825
rect 24766 36751 24822 36760
rect 25516 36145 25544 40967
rect 25608 40390 25636 41210
rect 25884 41206 25912 41482
rect 26146 41304 26202 41313
rect 26252 41274 26280 41618
rect 26146 41239 26202 41248
rect 26240 41268 26292 41274
rect 25872 41200 25924 41206
rect 25872 41142 25924 41148
rect 25962 40760 26018 40769
rect 25962 40695 26018 40704
rect 25596 40384 25648 40390
rect 25596 40326 25648 40332
rect 25608 39642 25636 40326
rect 25596 39636 25648 39642
rect 25596 39578 25648 39584
rect 25976 39409 26004 40695
rect 26160 40458 26188 41239
rect 26240 41210 26292 41216
rect 26240 40724 26292 40730
rect 26240 40666 26292 40672
rect 26148 40452 26200 40458
rect 26148 40394 26200 40400
rect 26056 39840 26108 39846
rect 26056 39782 26108 39788
rect 26068 39574 26096 39782
rect 26252 39642 26280 40666
rect 26344 40526 26372 42078
rect 26712 41750 26740 42502
rect 26896 42226 26924 43930
rect 27356 43926 27384 44134
rect 27344 43920 27396 43926
rect 27344 43862 27396 43868
rect 27068 43784 27120 43790
rect 27068 43726 27120 43732
rect 27080 42650 27108 43726
rect 27448 43296 27476 44270
rect 27724 43926 27752 44814
rect 28632 44328 28684 44334
rect 28632 44270 28684 44276
rect 27712 43920 27764 43926
rect 27712 43862 27764 43868
rect 28644 43450 28672 44270
rect 28724 44192 28776 44198
rect 28724 44134 28776 44140
rect 28632 43444 28684 43450
rect 28632 43386 28684 43392
rect 28264 43376 28316 43382
rect 28264 43318 28316 43324
rect 27620 43308 27672 43314
rect 27448 43268 27620 43296
rect 27252 43172 27304 43178
rect 27252 43114 27304 43120
rect 27264 42838 27292 43114
rect 27448 43110 27476 43268
rect 27620 43250 27672 43256
rect 27344 43104 27396 43110
rect 27344 43046 27396 43052
rect 27436 43104 27488 43110
rect 27436 43046 27488 43052
rect 27356 42838 27384 43046
rect 27252 42832 27304 42838
rect 27252 42774 27304 42780
rect 27344 42832 27396 42838
rect 27344 42774 27396 42780
rect 26988 42622 27108 42650
rect 26884 42220 26936 42226
rect 26884 42162 26936 42168
rect 26700 41744 26752 41750
rect 26700 41686 26752 41692
rect 26896 41138 26924 42162
rect 26988 41274 27016 42622
rect 27066 41984 27122 41993
rect 27066 41919 27122 41928
rect 27080 41818 27108 41919
rect 27068 41812 27120 41818
rect 27068 41754 27120 41760
rect 26976 41268 27028 41274
rect 26976 41210 27028 41216
rect 26884 41132 26936 41138
rect 26884 41074 26936 41080
rect 26424 40588 26476 40594
rect 26424 40530 26476 40536
rect 26516 40588 26568 40594
rect 26516 40530 26568 40536
rect 26332 40520 26384 40526
rect 26332 40462 26384 40468
rect 26436 39642 26464 40530
rect 26528 40186 26556 40530
rect 26792 40520 26844 40526
rect 26792 40462 26844 40468
rect 26884 40520 26936 40526
rect 26884 40462 26936 40468
rect 26700 40384 26752 40390
rect 26700 40326 26752 40332
rect 26712 40186 26740 40326
rect 26516 40180 26568 40186
rect 26516 40122 26568 40128
rect 26700 40180 26752 40186
rect 26700 40122 26752 40128
rect 26148 39636 26200 39642
rect 26148 39578 26200 39584
rect 26240 39636 26292 39642
rect 26240 39578 26292 39584
rect 26424 39636 26476 39642
rect 26424 39578 26476 39584
rect 26516 39636 26568 39642
rect 26516 39578 26568 39584
rect 26056 39568 26108 39574
rect 26056 39510 26108 39516
rect 26160 39438 26188 39578
rect 26240 39500 26292 39506
rect 26240 39442 26292 39448
rect 26148 39432 26200 39438
rect 25962 39400 26018 39409
rect 26148 39374 26200 39380
rect 25962 39335 26018 39344
rect 26252 38962 26280 39442
rect 26528 39438 26556 39578
rect 26516 39432 26568 39438
rect 26516 39374 26568 39380
rect 26804 39370 26832 40462
rect 26792 39364 26844 39370
rect 26792 39306 26844 39312
rect 26240 38956 26292 38962
rect 26240 38898 26292 38904
rect 26148 38888 26200 38894
rect 26148 38830 26200 38836
rect 25688 38752 25740 38758
rect 25686 38720 25688 38729
rect 25740 38720 25742 38729
rect 25686 38655 25742 38664
rect 26160 38593 26188 38830
rect 26146 38584 26202 38593
rect 26056 38548 26108 38554
rect 26146 38519 26202 38528
rect 26056 38490 26108 38496
rect 25688 38208 25740 38214
rect 25688 38150 25740 38156
rect 25700 38010 25728 38150
rect 25688 38004 25740 38010
rect 25688 37946 25740 37952
rect 26068 37097 26096 38490
rect 26148 38344 26200 38350
rect 26148 38286 26200 38292
rect 26160 37874 26188 38286
rect 26252 38282 26280 38898
rect 26804 38282 26832 39306
rect 26896 39030 26924 40462
rect 26988 40118 27016 41210
rect 27080 41070 27108 41754
rect 27448 41414 27476 43046
rect 27712 42900 27764 42906
rect 27712 42842 27764 42848
rect 27620 42696 27672 42702
rect 27620 42638 27672 42644
rect 27632 42226 27660 42638
rect 27620 42220 27672 42226
rect 27620 42162 27672 42168
rect 27724 41993 27752 42842
rect 28172 42696 28224 42702
rect 27802 42664 27858 42673
rect 28172 42638 28224 42644
rect 27802 42599 27804 42608
rect 27856 42599 27858 42608
rect 27804 42570 27856 42576
rect 27710 41984 27766 41993
rect 27710 41919 27766 41928
rect 28184 41818 28212 42638
rect 28276 42158 28304 43318
rect 28356 43308 28408 43314
rect 28356 43250 28408 43256
rect 28368 42702 28396 43250
rect 28736 43246 28764 44134
rect 28448 43240 28500 43246
rect 28448 43182 28500 43188
rect 28724 43240 28776 43246
rect 28724 43182 28776 43188
rect 28356 42696 28408 42702
rect 28356 42638 28408 42644
rect 28264 42152 28316 42158
rect 28264 42094 28316 42100
rect 27528 41812 27580 41818
rect 27528 41754 27580 41760
rect 28172 41812 28224 41818
rect 28172 41754 28224 41760
rect 27264 41386 27476 41414
rect 27160 41268 27212 41274
rect 27160 41210 27212 41216
rect 27172 41177 27200 41210
rect 27158 41168 27214 41177
rect 27158 41103 27214 41112
rect 27068 41064 27120 41070
rect 27068 41006 27120 41012
rect 27066 40624 27122 40633
rect 27066 40559 27122 40568
rect 27080 40526 27108 40559
rect 27068 40520 27120 40526
rect 27068 40462 27120 40468
rect 26976 40112 27028 40118
rect 26976 40054 27028 40060
rect 26976 39636 27028 39642
rect 26976 39578 27028 39584
rect 26884 39024 26936 39030
rect 26884 38966 26936 38972
rect 26884 38344 26936 38350
rect 26884 38286 26936 38292
rect 26240 38276 26292 38282
rect 26240 38218 26292 38224
rect 26792 38276 26844 38282
rect 26792 38218 26844 38224
rect 26148 37868 26200 37874
rect 26148 37810 26200 37816
rect 26252 37262 26280 38218
rect 26896 38010 26924 38286
rect 26884 38004 26936 38010
rect 26884 37946 26936 37952
rect 26516 37732 26568 37738
rect 26516 37674 26568 37680
rect 26528 37466 26556 37674
rect 26516 37460 26568 37466
rect 26516 37402 26568 37408
rect 26240 37256 26292 37262
rect 26240 37198 26292 37204
rect 26054 37088 26110 37097
rect 26054 37023 26110 37032
rect 25872 36848 25924 36854
rect 25872 36790 25924 36796
rect 25502 36136 25558 36145
rect 24492 36100 24544 36106
rect 25502 36071 25558 36080
rect 24492 36042 24544 36048
rect 24308 35964 24360 35970
rect 24308 35906 24360 35912
rect 24504 35873 24532 36042
rect 25228 36032 25280 36038
rect 25228 35974 25280 35980
rect 24768 35896 24820 35902
rect 23570 35864 23626 35873
rect 23570 35799 23626 35808
rect 24490 35864 24546 35873
rect 24490 35799 24546 35808
rect 24766 35864 24768 35873
rect 24820 35864 24822 35873
rect 24766 35799 24822 35808
rect 25240 35737 25268 35974
rect 25884 35873 25912 36790
rect 26988 36514 27016 39578
rect 27264 39506 27292 41386
rect 27436 41064 27488 41070
rect 27436 41006 27488 41012
rect 27344 39908 27396 39914
rect 27344 39850 27396 39856
rect 27356 39642 27384 39850
rect 27448 39846 27476 41006
rect 27540 40934 27568 41754
rect 27712 41540 27764 41546
rect 27712 41482 27764 41488
rect 27724 41449 27752 41482
rect 27710 41440 27766 41449
rect 28276 41414 28304 42094
rect 28460 41614 28488 43182
rect 28632 43172 28684 43178
rect 28632 43114 28684 43120
rect 28644 42702 28672 43114
rect 28828 42770 28856 44814
rect 29184 44736 29236 44742
rect 29184 44678 29236 44684
rect 29196 44266 29224 44678
rect 30944 44538 30972 44814
rect 31758 44775 31814 44784
rect 33508 44804 33560 44810
rect 30932 44532 30984 44538
rect 30932 44474 30984 44480
rect 30472 44328 30524 44334
rect 30472 44270 30524 44276
rect 29184 44260 29236 44266
rect 29184 44202 29236 44208
rect 28908 43852 28960 43858
rect 28908 43794 28960 43800
rect 28920 43382 28948 43794
rect 29000 43784 29052 43790
rect 29000 43726 29052 43732
rect 29012 43450 29040 43726
rect 29000 43444 29052 43450
rect 29000 43386 29052 43392
rect 28908 43376 28960 43382
rect 28908 43318 28960 43324
rect 29092 43104 29144 43110
rect 29092 43046 29144 43052
rect 29000 42832 29052 42838
rect 29000 42774 29052 42780
rect 28816 42764 28868 42770
rect 28816 42706 28868 42712
rect 28632 42696 28684 42702
rect 28632 42638 28684 42644
rect 28644 42362 28672 42638
rect 29012 42362 29040 42774
rect 29104 42702 29132 43046
rect 29092 42696 29144 42702
rect 29092 42638 29144 42644
rect 28632 42356 28684 42362
rect 28632 42298 28684 42304
rect 29000 42356 29052 42362
rect 29000 42298 29052 42304
rect 28540 42288 28592 42294
rect 28540 42230 28592 42236
rect 28552 41682 28580 42230
rect 28644 42158 28672 42298
rect 28632 42152 28684 42158
rect 28632 42094 28684 42100
rect 28722 41848 28778 41857
rect 28722 41783 28778 41792
rect 28540 41676 28592 41682
rect 28540 41618 28592 41624
rect 28448 41608 28500 41614
rect 28448 41550 28500 41556
rect 28552 41414 28580 41618
rect 27710 41375 27766 41384
rect 28000 41386 28304 41414
rect 28460 41386 28580 41414
rect 27528 40928 27580 40934
rect 27528 40870 27580 40876
rect 27528 40520 27580 40526
rect 27528 40462 27580 40468
rect 27436 39840 27488 39846
rect 27436 39782 27488 39788
rect 27344 39636 27396 39642
rect 27344 39578 27396 39584
rect 27448 39506 27476 39782
rect 27252 39500 27304 39506
rect 27252 39442 27304 39448
rect 27436 39500 27488 39506
rect 27436 39442 27488 39448
rect 27540 39386 27568 40462
rect 27710 40352 27766 40361
rect 27710 40287 27766 40296
rect 27620 39568 27672 39574
rect 27620 39510 27672 39516
rect 27448 39358 27568 39386
rect 27448 37262 27476 39358
rect 27632 38894 27660 39510
rect 27620 38888 27672 38894
rect 27620 38830 27672 38836
rect 27724 38706 27752 40287
rect 28000 40186 28028 41386
rect 28080 40384 28132 40390
rect 28080 40326 28132 40332
rect 27988 40180 28040 40186
rect 27988 40122 28040 40128
rect 27802 38856 27858 38865
rect 27802 38791 27804 38800
rect 27856 38791 27858 38800
rect 27804 38762 27856 38768
rect 27540 38678 27752 38706
rect 27540 38554 27568 38678
rect 27528 38548 27580 38554
rect 27528 38490 27580 38496
rect 27620 38548 27672 38554
rect 27620 38490 27672 38496
rect 27632 38457 27660 38490
rect 27618 38448 27674 38457
rect 27618 38383 27674 38392
rect 27804 38344 27856 38350
rect 27804 38286 27856 38292
rect 27620 37936 27672 37942
rect 27620 37878 27672 37884
rect 27632 37806 27660 37878
rect 27620 37800 27672 37806
rect 27620 37742 27672 37748
rect 27816 37670 27844 38286
rect 28000 37942 28028 40122
rect 28092 39642 28120 40326
rect 28460 40066 28488 41386
rect 28460 40038 28672 40066
rect 28644 39914 28672 40038
rect 28632 39908 28684 39914
rect 28632 39850 28684 39856
rect 28080 39636 28132 39642
rect 28080 39578 28132 39584
rect 28172 39432 28224 39438
rect 28172 39374 28224 39380
rect 28184 38282 28212 39374
rect 28540 38888 28592 38894
rect 28540 38830 28592 38836
rect 28172 38276 28224 38282
rect 28172 38218 28224 38224
rect 27988 37936 28040 37942
rect 27988 37878 28040 37884
rect 27896 37800 27948 37806
rect 27896 37742 27948 37748
rect 27804 37664 27856 37670
rect 27804 37606 27856 37612
rect 27816 37466 27844 37606
rect 27804 37460 27856 37466
rect 27804 37402 27856 37408
rect 27908 37369 27936 37742
rect 28552 37670 28580 38830
rect 28644 38826 28672 39850
rect 28632 38820 28684 38826
rect 28632 38762 28684 38768
rect 28632 38208 28684 38214
rect 28632 38150 28684 38156
rect 28644 37874 28672 38150
rect 28632 37868 28684 37874
rect 28632 37810 28684 37816
rect 28540 37664 28592 37670
rect 28540 37606 28592 37612
rect 28552 37369 28580 37606
rect 27894 37360 27950 37369
rect 27894 37295 27950 37304
rect 28538 37360 28594 37369
rect 28538 37295 28594 37304
rect 27436 37256 27488 37262
rect 27436 37198 27488 37204
rect 27620 37120 27672 37126
rect 27620 37062 27672 37068
rect 26976 36508 27028 36514
rect 26976 36450 27028 36456
rect 25870 35864 25926 35873
rect 27632 35834 27660 37062
rect 28736 36242 28764 41783
rect 29104 41596 29132 42638
rect 29196 42634 29224 44202
rect 29368 44192 29420 44198
rect 29368 44134 29420 44140
rect 29380 43246 29408 44134
rect 29644 43920 29696 43926
rect 29644 43862 29696 43868
rect 29656 43450 29684 43862
rect 30380 43784 30432 43790
rect 30484 43738 30512 44270
rect 30840 44260 30892 44266
rect 30840 44202 30892 44208
rect 30748 44192 30800 44198
rect 30748 44134 30800 44140
rect 30656 43852 30708 43858
rect 30656 43794 30708 43800
rect 30432 43732 30512 43738
rect 30380 43726 30512 43732
rect 30392 43710 30512 43726
rect 29644 43444 29696 43450
rect 29644 43386 29696 43392
rect 30104 43444 30156 43450
rect 30104 43386 30156 43392
rect 29642 43344 29698 43353
rect 30116 43314 30144 43386
rect 29642 43279 29644 43288
rect 29696 43279 29698 43288
rect 30104 43308 30156 43314
rect 29644 43250 29696 43256
rect 30104 43250 30156 43256
rect 29368 43240 29420 43246
rect 29368 43182 29420 43188
rect 29736 43104 29788 43110
rect 29736 43046 29788 43052
rect 29748 42634 29776 43046
rect 29184 42628 29236 42634
rect 29184 42570 29236 42576
rect 29736 42628 29788 42634
rect 29736 42570 29788 42576
rect 30116 42566 30144 43250
rect 30196 43172 30248 43178
rect 30196 43114 30248 43120
rect 30208 42838 30236 43114
rect 30288 43104 30340 43110
rect 30288 43046 30340 43052
rect 30196 42832 30248 42838
rect 30196 42774 30248 42780
rect 30300 42634 30328 43046
rect 30380 42832 30432 42838
rect 30380 42774 30432 42780
rect 30288 42628 30340 42634
rect 30288 42570 30340 42576
rect 30104 42560 30156 42566
rect 30104 42502 30156 42508
rect 30116 41682 30144 42502
rect 30196 42152 30248 42158
rect 30196 42094 30248 42100
rect 30104 41676 30156 41682
rect 30104 41618 30156 41624
rect 29184 41608 29236 41614
rect 29104 41568 29184 41596
rect 29184 41550 29236 41556
rect 30104 41064 30156 41070
rect 30104 41006 30156 41012
rect 29092 40928 29144 40934
rect 29092 40870 29144 40876
rect 29920 40928 29972 40934
rect 29920 40870 29972 40876
rect 29104 40730 29132 40870
rect 29092 40724 29144 40730
rect 29092 40666 29144 40672
rect 29932 40662 29960 40870
rect 29920 40656 29972 40662
rect 29920 40598 29972 40604
rect 30012 40656 30064 40662
rect 30012 40598 30064 40604
rect 28816 40588 28868 40594
rect 28816 40530 28868 40536
rect 28828 40186 28856 40530
rect 29276 40520 29328 40526
rect 29274 40488 29276 40497
rect 29368 40520 29420 40526
rect 29328 40488 29330 40497
rect 29368 40462 29420 40468
rect 29274 40423 29330 40432
rect 29276 40384 29328 40390
rect 29276 40326 29328 40332
rect 28816 40180 28868 40186
rect 28816 40122 28868 40128
rect 28908 39840 28960 39846
rect 28908 39782 28960 39788
rect 28814 39672 28870 39681
rect 28814 39607 28870 39616
rect 28828 39438 28856 39607
rect 28920 39574 28948 39782
rect 28908 39568 28960 39574
rect 29090 39536 29146 39545
rect 28908 39510 28960 39516
rect 29012 39494 29090 39522
rect 28816 39432 28868 39438
rect 28816 39374 28868 39380
rect 29012 39250 29040 39494
rect 29090 39471 29146 39480
rect 28966 39222 29040 39250
rect 28966 39098 28994 39222
rect 29288 39098 29316 40326
rect 29380 40050 29408 40462
rect 29734 40216 29790 40225
rect 29734 40151 29790 40160
rect 29368 40044 29420 40050
rect 29368 39986 29420 39992
rect 29380 39386 29408 39986
rect 29748 39642 29776 40151
rect 29828 39908 29880 39914
rect 29828 39850 29880 39856
rect 29736 39636 29788 39642
rect 29736 39578 29788 39584
rect 29642 39536 29698 39545
rect 29642 39471 29698 39480
rect 29380 39358 29592 39386
rect 29380 39302 29408 39358
rect 29368 39296 29420 39302
rect 29368 39238 29420 39244
rect 29460 39296 29512 39302
rect 29460 39238 29512 39244
rect 28954 39092 29006 39098
rect 28954 39034 29006 39040
rect 29276 39092 29328 39098
rect 29276 39034 29328 39040
rect 28908 38956 28960 38962
rect 28960 38916 29224 38944
rect 28908 38898 28960 38904
rect 28954 38752 29006 38758
rect 29092 38752 29144 38758
rect 29006 38712 29092 38740
rect 28954 38694 29006 38700
rect 29092 38694 29144 38700
rect 29196 38654 29224 38916
rect 29472 38865 29500 39238
rect 29458 38856 29514 38865
rect 29458 38791 29514 38800
rect 29564 38654 29592 39358
rect 29656 39098 29684 39471
rect 29644 39092 29696 39098
rect 29644 39034 29696 39040
rect 29104 38626 29224 38654
rect 29380 38626 29592 38654
rect 29000 37392 29052 37398
rect 29000 37334 29052 37340
rect 28816 36508 28868 36514
rect 28816 36450 28868 36456
rect 28828 36242 28856 36450
rect 29012 36281 29040 37334
rect 29104 37097 29132 38626
rect 29184 38344 29236 38350
rect 29184 38286 29236 38292
rect 29196 37738 29224 38286
rect 29184 37732 29236 37738
rect 29184 37674 29236 37680
rect 29196 37466 29224 37674
rect 29184 37460 29236 37466
rect 29184 37402 29236 37408
rect 29380 37330 29408 38626
rect 29840 38486 29868 39850
rect 29920 39500 29972 39506
rect 30024 39488 30052 40598
rect 30116 40050 30144 41006
rect 30104 40044 30156 40050
rect 30104 39986 30156 39992
rect 30116 39574 30144 39986
rect 30104 39568 30156 39574
rect 30104 39510 30156 39516
rect 29972 39460 30052 39488
rect 29920 39442 29972 39448
rect 30012 38956 30064 38962
rect 30116 38944 30144 39510
rect 30064 38916 30144 38944
rect 30012 38898 30064 38904
rect 29828 38480 29880 38486
rect 29828 38422 29880 38428
rect 30012 38344 30064 38350
rect 29550 38312 29606 38321
rect 30012 38286 30064 38292
rect 29550 38247 29552 38256
rect 29604 38247 29606 38256
rect 29552 38218 29604 38224
rect 30024 37670 30052 38286
rect 29644 37664 29696 37670
rect 29644 37606 29696 37612
rect 30012 37664 30064 37670
rect 30012 37606 30064 37612
rect 29656 37398 29684 37606
rect 29920 37460 29972 37466
rect 29920 37402 29972 37408
rect 29644 37392 29696 37398
rect 29644 37334 29696 37340
rect 29368 37324 29420 37330
rect 29368 37266 29420 37272
rect 29090 37088 29146 37097
rect 29090 37023 29146 37032
rect 28998 36272 29054 36281
rect 28724 36236 28776 36242
rect 28724 36178 28776 36184
rect 28816 36236 28868 36242
rect 28998 36207 29054 36216
rect 28816 36178 28868 36184
rect 25870 35799 25926 35808
rect 27620 35828 27672 35834
rect 27620 35770 27672 35776
rect 14832 35702 14884 35708
rect 15014 35728 15070 35737
rect 8206 35663 8262 35672
rect 15014 35663 15070 35672
rect 20074 35728 20130 35737
rect 20074 35663 20130 35672
rect 21362 35728 21418 35737
rect 21362 35663 21418 35672
rect 22190 35728 22246 35737
rect 22190 35663 22192 35672
rect 22244 35663 22246 35672
rect 23018 35728 23074 35737
rect 23018 35663 23074 35672
rect 23202 35728 23258 35737
rect 23202 35663 23258 35672
rect 25226 35728 25282 35737
rect 25226 35663 25282 35672
rect 22192 35634 22244 35640
rect 23032 35630 23060 35663
rect 23020 35624 23072 35630
rect 23020 35566 23072 35572
rect 29932 35578 29960 37402
rect 30024 35873 30052 37606
rect 30102 36544 30158 36553
rect 30102 36479 30158 36488
rect 30116 35902 30144 36479
rect 30104 35896 30156 35902
rect 30010 35864 30066 35873
rect 30208 35873 30236 42094
rect 30392 42022 30420 42774
rect 30484 42770 30512 43710
rect 30562 43480 30618 43489
rect 30562 43415 30618 43424
rect 30576 43246 30604 43415
rect 30564 43240 30616 43246
rect 30564 43182 30616 43188
rect 30564 43104 30616 43110
rect 30668 43092 30696 43794
rect 30760 43382 30788 44134
rect 30748 43376 30800 43382
rect 30748 43318 30800 43324
rect 30616 43064 30696 43092
rect 30564 43046 30616 43052
rect 30472 42764 30524 42770
rect 30472 42706 30524 42712
rect 30380 42016 30432 42022
rect 30378 41984 30380 41993
rect 30472 42016 30524 42022
rect 30432 41984 30434 41993
rect 30472 41958 30524 41964
rect 30378 41919 30434 41928
rect 30380 41540 30432 41546
rect 30380 41482 30432 41488
rect 30392 41414 30420 41482
rect 30484 41478 30512 41958
rect 30472 41472 30524 41478
rect 30472 41414 30524 41420
rect 30300 41386 30420 41414
rect 30300 40186 30328 41386
rect 30378 41032 30434 41041
rect 30378 40967 30434 40976
rect 30392 40526 30420 40967
rect 30576 40730 30604 43046
rect 30760 42090 30788 43318
rect 30852 42294 30880 44202
rect 31392 43784 31444 43790
rect 31390 43752 31392 43761
rect 31444 43752 31446 43761
rect 31390 43687 31446 43696
rect 31206 43344 31262 43353
rect 31206 43279 31262 43288
rect 31220 43246 31248 43279
rect 31208 43240 31260 43246
rect 31208 43182 31260 43188
rect 31404 43178 31432 43687
rect 31668 43648 31720 43654
rect 31668 43590 31720 43596
rect 31680 43489 31708 43590
rect 31666 43480 31722 43489
rect 31576 43444 31628 43450
rect 31666 43415 31722 43424
rect 31576 43386 31628 43392
rect 31588 43246 31616 43386
rect 31576 43240 31628 43246
rect 31576 43182 31628 43188
rect 31392 43172 31444 43178
rect 31392 43114 31444 43120
rect 30840 42288 30892 42294
rect 30840 42230 30892 42236
rect 30656 42084 30708 42090
rect 30656 42026 30708 42032
rect 30748 42084 30800 42090
rect 30748 42026 30800 42032
rect 30668 41478 30696 42026
rect 31114 41984 31170 41993
rect 31114 41919 31170 41928
rect 30840 41744 30892 41750
rect 31128 41721 31156 41919
rect 30840 41686 30892 41692
rect 31114 41712 31170 41721
rect 30656 41472 30708 41478
rect 30656 41414 30708 41420
rect 30656 41064 30708 41070
rect 30656 41006 30708 41012
rect 30668 40730 30696 41006
rect 30564 40724 30616 40730
rect 30564 40666 30616 40672
rect 30656 40724 30708 40730
rect 30656 40666 30708 40672
rect 30380 40520 30432 40526
rect 30380 40462 30432 40468
rect 30472 40384 30524 40390
rect 30472 40326 30524 40332
rect 30484 40186 30512 40326
rect 30288 40180 30340 40186
rect 30288 40122 30340 40128
rect 30472 40180 30524 40186
rect 30472 40122 30524 40128
rect 30300 37874 30328 40122
rect 30576 40050 30604 40666
rect 30564 40044 30616 40050
rect 30564 39986 30616 39992
rect 30576 39914 30604 39986
rect 30380 39908 30432 39914
rect 30380 39850 30432 39856
rect 30564 39908 30616 39914
rect 30564 39850 30616 39856
rect 30392 39642 30420 39850
rect 30748 39840 30800 39846
rect 30748 39782 30800 39788
rect 30380 39636 30432 39642
rect 30380 39578 30432 39584
rect 30472 39500 30524 39506
rect 30472 39442 30524 39448
rect 30380 39364 30432 39370
rect 30484 39352 30512 39442
rect 30432 39324 30512 39352
rect 30380 39306 30432 39312
rect 30484 38418 30512 39324
rect 30564 38956 30616 38962
rect 30564 38898 30616 38904
rect 30576 38486 30604 38898
rect 30760 38740 30788 39782
rect 30852 39545 30880 41686
rect 31114 41647 31170 41656
rect 31576 41540 31628 41546
rect 31576 41482 31628 41488
rect 31588 41138 31616 41482
rect 31116 41132 31168 41138
rect 31116 41074 31168 41080
rect 31576 41132 31628 41138
rect 31576 41074 31628 41080
rect 30838 39536 30894 39545
rect 30838 39471 30894 39480
rect 30840 39432 30892 39438
rect 30840 39374 30892 39380
rect 30852 39030 30880 39374
rect 30840 39024 30892 39030
rect 30840 38966 30892 38972
rect 31128 38962 31156 41074
rect 31208 40520 31260 40526
rect 31206 40488 31208 40497
rect 31260 40488 31262 40497
rect 31206 40423 31262 40432
rect 31220 39438 31248 40423
rect 31588 40118 31616 41074
rect 31666 40624 31722 40633
rect 31666 40559 31668 40568
rect 31720 40559 31722 40568
rect 31668 40530 31720 40536
rect 31576 40112 31628 40118
rect 31576 40054 31628 40060
rect 31300 40044 31352 40050
rect 31300 39986 31352 39992
rect 31392 40044 31444 40050
rect 31392 39986 31444 39992
rect 31312 39642 31340 39986
rect 31300 39636 31352 39642
rect 31300 39578 31352 39584
rect 31208 39432 31260 39438
rect 31208 39374 31260 39380
rect 31404 39302 31432 39986
rect 31576 39840 31628 39846
rect 31576 39782 31628 39788
rect 31392 39296 31444 39302
rect 31392 39238 31444 39244
rect 31116 38956 31168 38962
rect 31116 38898 31168 38904
rect 30840 38752 30892 38758
rect 30760 38712 30840 38740
rect 30840 38694 30892 38700
rect 30564 38480 30616 38486
rect 30564 38422 30616 38428
rect 30748 38480 30800 38486
rect 30748 38422 30800 38428
rect 30472 38412 30524 38418
rect 30472 38354 30524 38360
rect 30656 38208 30708 38214
rect 30656 38150 30708 38156
rect 30668 37942 30696 38150
rect 30656 37936 30708 37942
rect 30656 37878 30708 37884
rect 30288 37868 30340 37874
rect 30288 37810 30340 37816
rect 30656 37800 30708 37806
rect 30760 37754 30788 38422
rect 31128 38350 31156 38898
rect 31588 38826 31616 39782
rect 31576 38820 31628 38826
rect 31576 38762 31628 38768
rect 31208 38752 31260 38758
rect 31206 38720 31208 38729
rect 31392 38752 31444 38758
rect 31260 38720 31262 38729
rect 31392 38694 31444 38700
rect 31206 38655 31262 38664
rect 31404 38418 31432 38694
rect 31392 38412 31444 38418
rect 31392 38354 31444 38360
rect 31116 38344 31168 38350
rect 31116 38286 31168 38292
rect 31484 38344 31536 38350
rect 31484 38286 31536 38292
rect 30708 37748 30788 37754
rect 30656 37742 30788 37748
rect 30668 37726 30788 37742
rect 30668 37398 30696 37726
rect 30656 37392 30708 37398
rect 30656 37334 30708 37340
rect 30378 36816 30434 36825
rect 30378 36751 30434 36760
rect 30288 36576 30340 36582
rect 30288 36518 30340 36524
rect 30104 35838 30156 35844
rect 30194 35864 30250 35873
rect 30010 35799 30066 35808
rect 30194 35799 30250 35808
rect 30300 35737 30328 36518
rect 30392 36514 30420 36751
rect 30472 36644 30524 36650
rect 30472 36586 30524 36592
rect 30380 36508 30432 36514
rect 30380 36450 30432 36456
rect 30484 36417 30512 36586
rect 30470 36408 30526 36417
rect 30470 36343 30526 36352
rect 31128 35873 31156 38286
rect 31496 37126 31524 38286
rect 31668 37732 31720 37738
rect 31668 37674 31720 37680
rect 31680 37466 31708 37674
rect 31668 37460 31720 37466
rect 31668 37402 31720 37408
rect 31772 37398 31800 44775
rect 33508 44746 33560 44752
rect 33048 44396 33100 44402
rect 33048 44338 33100 44344
rect 31852 44328 31904 44334
rect 31852 44270 31904 44276
rect 31864 43858 31892 44270
rect 32404 44192 32456 44198
rect 32404 44134 32456 44140
rect 31852 43852 31904 43858
rect 31852 43794 31904 43800
rect 32220 43784 32272 43790
rect 32220 43726 32272 43732
rect 32128 43716 32180 43722
rect 32128 43658 32180 43664
rect 32140 42702 32168 43658
rect 32232 43110 32260 43726
rect 32220 43104 32272 43110
rect 32220 43046 32272 43052
rect 32416 42838 32444 44134
rect 33060 43790 33088 44338
rect 33324 44192 33376 44198
rect 33324 44134 33376 44140
rect 33416 44192 33468 44198
rect 33416 44134 33468 44140
rect 33048 43784 33100 43790
rect 33048 43726 33100 43732
rect 33232 43648 33284 43654
rect 33232 43590 33284 43596
rect 33140 43444 33192 43450
rect 33140 43386 33192 43392
rect 32404 42832 32456 42838
rect 32404 42774 32456 42780
rect 32128 42696 32180 42702
rect 31850 42664 31906 42673
rect 32128 42638 32180 42644
rect 31850 42599 31906 42608
rect 31864 42090 31892 42599
rect 31852 42084 31904 42090
rect 31852 42026 31904 42032
rect 31944 41608 31996 41614
rect 31850 41576 31906 41585
rect 31944 41550 31996 41556
rect 31850 41511 31852 41520
rect 31904 41511 31906 41520
rect 31852 41482 31904 41488
rect 31850 41032 31906 41041
rect 31850 40967 31852 40976
rect 31904 40967 31906 40976
rect 31852 40938 31904 40944
rect 31852 40520 31904 40526
rect 31852 40462 31904 40468
rect 31864 40390 31892 40462
rect 31852 40384 31904 40390
rect 31852 40326 31904 40332
rect 31864 39284 31892 40326
rect 31956 39506 31984 41550
rect 32036 41472 32088 41478
rect 32036 41414 32088 41420
rect 32048 40089 32076 41414
rect 32140 41138 32168 42638
rect 32494 42528 32550 42537
rect 32494 42463 32550 42472
rect 32312 42220 32364 42226
rect 32312 42162 32364 42168
rect 32220 42016 32272 42022
rect 32220 41958 32272 41964
rect 32232 41750 32260 41958
rect 32220 41744 32272 41750
rect 32220 41686 32272 41692
rect 32128 41132 32180 41138
rect 32324 41120 32352 42162
rect 32404 42084 32456 42090
rect 32404 42026 32456 42032
rect 32416 41478 32444 42026
rect 32404 41472 32456 41478
rect 32404 41414 32456 41420
rect 32324 41092 32444 41120
rect 32128 41074 32180 41080
rect 32140 40662 32168 41074
rect 32220 40928 32272 40934
rect 32220 40870 32272 40876
rect 32128 40656 32180 40662
rect 32128 40598 32180 40604
rect 32128 40384 32180 40390
rect 32128 40326 32180 40332
rect 32034 40080 32090 40089
rect 32034 40015 32090 40024
rect 32140 39574 32168 40326
rect 32128 39568 32180 39574
rect 32128 39510 32180 39516
rect 31944 39500 31996 39506
rect 31996 39460 32076 39488
rect 31944 39442 31996 39448
rect 31864 39256 31984 39284
rect 31956 37754 31984 39256
rect 32048 37874 32076 39460
rect 32232 39030 32260 40870
rect 32220 39024 32272 39030
rect 32220 38966 32272 38972
rect 32128 38956 32180 38962
rect 32128 38898 32180 38904
rect 32140 38758 32168 38898
rect 32128 38752 32180 38758
rect 32128 38694 32180 38700
rect 32220 38208 32272 38214
rect 32220 38150 32272 38156
rect 32036 37868 32088 37874
rect 32036 37810 32088 37816
rect 31852 37732 31904 37738
rect 31956 37726 32076 37754
rect 31852 37674 31904 37680
rect 31864 37466 31892 37674
rect 31852 37460 31904 37466
rect 31852 37402 31904 37408
rect 31760 37392 31812 37398
rect 31760 37334 31812 37340
rect 31864 37330 31892 37402
rect 31852 37324 31904 37330
rect 31852 37266 31904 37272
rect 31944 37324 31996 37330
rect 31944 37266 31996 37272
rect 31484 37120 31536 37126
rect 31484 37062 31536 37068
rect 31956 36922 31984 37266
rect 32048 37262 32076 37726
rect 32232 37466 32260 38150
rect 32220 37460 32272 37466
rect 32220 37402 32272 37408
rect 32036 37256 32088 37262
rect 32416 37233 32444 41092
rect 32508 39386 32536 42463
rect 33046 42256 33102 42265
rect 33152 42226 33180 43386
rect 33244 43178 33272 43590
rect 33336 43450 33364 44134
rect 33324 43444 33376 43450
rect 33324 43386 33376 43392
rect 33232 43172 33284 43178
rect 33232 43114 33284 43120
rect 33428 42634 33456 44134
rect 33416 42628 33468 42634
rect 33416 42570 33468 42576
rect 33520 42265 33548 44746
rect 34244 44328 34296 44334
rect 34244 44270 34296 44276
rect 33968 44192 34020 44198
rect 33968 44134 34020 44140
rect 33980 43926 34008 44134
rect 33968 43920 34020 43926
rect 33968 43862 34020 43868
rect 34060 43920 34112 43926
rect 34060 43862 34112 43868
rect 33600 43784 33652 43790
rect 33600 43726 33652 43732
rect 33612 42362 33640 43726
rect 33692 43648 33744 43654
rect 33692 43590 33744 43596
rect 33704 43314 33732 43590
rect 33692 43308 33744 43314
rect 33692 43250 33744 43256
rect 34072 43178 34100 43862
rect 34256 43450 34284 44270
rect 34336 43648 34388 43654
rect 34336 43590 34388 43596
rect 34244 43444 34296 43450
rect 34244 43386 34296 43392
rect 33692 43172 33744 43178
rect 33692 43114 33744 43120
rect 34060 43172 34112 43178
rect 34060 43114 34112 43120
rect 33704 42838 33732 43114
rect 33692 42832 33744 42838
rect 33692 42774 33744 42780
rect 33692 42696 33744 42702
rect 33692 42638 33744 42644
rect 33600 42356 33652 42362
rect 33600 42298 33652 42304
rect 33506 42256 33562 42265
rect 33046 42191 33102 42200
rect 33140 42220 33192 42226
rect 33060 42106 33088 42191
rect 33140 42162 33192 42168
rect 33416 42220 33468 42226
rect 33506 42191 33562 42200
rect 33416 42162 33468 42168
rect 33060 42078 33364 42106
rect 33428 42090 33456 42162
rect 33704 42158 33732 42638
rect 33692 42152 33744 42158
rect 33692 42094 33744 42100
rect 33336 42022 33364 42078
rect 33416 42084 33468 42090
rect 33416 42026 33468 42032
rect 33232 42016 33284 42022
rect 33232 41958 33284 41964
rect 33324 42016 33376 42022
rect 33324 41958 33376 41964
rect 33244 40730 33272 41958
rect 33704 41818 33732 42094
rect 33692 41812 33744 41818
rect 33692 41754 33744 41760
rect 33324 41676 33376 41682
rect 33324 41618 33376 41624
rect 33232 40724 33284 40730
rect 33232 40666 33284 40672
rect 33048 40656 33100 40662
rect 33048 40598 33100 40604
rect 32956 40520 33008 40526
rect 32956 40462 33008 40468
rect 32588 39908 32640 39914
rect 32588 39850 32640 39856
rect 32600 39642 32628 39850
rect 32968 39846 32996 40462
rect 32956 39840 33008 39846
rect 32862 39808 32918 39817
rect 32956 39782 33008 39788
rect 32862 39743 32918 39752
rect 32588 39636 32640 39642
rect 32588 39578 32640 39584
rect 32508 39358 32628 39386
rect 32494 39264 32550 39273
rect 32494 39199 32550 39208
rect 32508 38865 32536 39199
rect 32494 38856 32550 38865
rect 32494 38791 32550 38800
rect 32600 37466 32628 39358
rect 32680 39296 32732 39302
rect 32678 39264 32680 39273
rect 32772 39296 32824 39302
rect 32732 39264 32734 39273
rect 32772 39238 32824 39244
rect 32678 39199 32734 39208
rect 32784 39137 32812 39238
rect 32770 39128 32826 39137
rect 32770 39063 32826 39072
rect 32784 38826 32812 39063
rect 32772 38820 32824 38826
rect 32772 38762 32824 38768
rect 32588 37460 32640 37466
rect 32588 37402 32640 37408
rect 32036 37198 32088 37204
rect 32402 37224 32458 37233
rect 32402 37159 32458 37168
rect 31668 36916 31720 36922
rect 31668 36858 31720 36864
rect 31944 36916 31996 36922
rect 31944 36858 31996 36864
rect 31680 36009 31708 36858
rect 32876 36417 32904 39743
rect 32968 39409 32996 39782
rect 32954 39400 33010 39409
rect 32954 39335 33010 39344
rect 33060 38434 33088 40598
rect 33140 40588 33192 40594
rect 33140 40530 33192 40536
rect 33152 39642 33180 40530
rect 33336 39914 33364 41618
rect 33508 41540 33560 41546
rect 33508 41482 33560 41488
rect 33416 40928 33468 40934
rect 33416 40870 33468 40876
rect 33324 39908 33376 39914
rect 33324 39850 33376 39856
rect 33140 39636 33192 39642
rect 33140 39578 33192 39584
rect 33060 38418 33180 38434
rect 33060 38412 33192 38418
rect 33060 38406 33140 38412
rect 33140 38354 33192 38360
rect 33138 37904 33194 37913
rect 33060 37862 33138 37890
rect 33060 36446 33088 37862
rect 33138 37839 33194 37848
rect 33048 36440 33100 36446
rect 32862 36408 32918 36417
rect 33048 36382 33100 36388
rect 32862 36343 32918 36352
rect 33048 36236 33100 36242
rect 33048 36178 33100 36184
rect 31666 36000 31722 36009
rect 31666 35935 31722 35944
rect 33060 35873 33088 36178
rect 33428 36009 33456 40870
rect 33520 40526 33548 41482
rect 33704 40730 33732 41754
rect 34072 41682 34100 43114
rect 34348 43110 34376 43590
rect 34612 43240 34664 43246
rect 34612 43182 34664 43188
rect 34336 43104 34388 43110
rect 34336 43046 34388 43052
rect 34348 42838 34376 43046
rect 34152 42832 34204 42838
rect 34152 42774 34204 42780
rect 34336 42832 34388 42838
rect 34336 42774 34388 42780
rect 34060 41676 34112 41682
rect 34060 41618 34112 41624
rect 33876 41608 33928 41614
rect 33876 41550 33928 41556
rect 33888 41274 33916 41550
rect 33876 41268 33928 41274
rect 33876 41210 33928 41216
rect 33692 40724 33744 40730
rect 33692 40666 33744 40672
rect 33784 40588 33836 40594
rect 33888 40576 33916 41210
rect 34164 41002 34192 42774
rect 34520 42696 34572 42702
rect 34440 42644 34520 42650
rect 34440 42638 34572 42644
rect 34440 42622 34560 42638
rect 34440 42158 34468 42622
rect 34624 42566 34652 43182
rect 35164 43172 35216 43178
rect 35164 43114 35216 43120
rect 35072 42764 35124 42770
rect 35072 42706 35124 42712
rect 34980 42696 35032 42702
rect 34980 42638 35032 42644
rect 34612 42560 34664 42566
rect 34612 42502 34664 42508
rect 34624 42226 34652 42502
rect 34796 42288 34848 42294
rect 34796 42230 34848 42236
rect 34612 42220 34664 42226
rect 34612 42162 34664 42168
rect 34428 42152 34480 42158
rect 34428 42094 34480 42100
rect 34244 42084 34296 42090
rect 34244 42026 34296 42032
rect 34256 41138 34284 42026
rect 34440 41546 34468 42094
rect 34428 41540 34480 41546
rect 34428 41482 34480 41488
rect 34520 41472 34572 41478
rect 34518 41440 34520 41449
rect 34572 41440 34574 41449
rect 34518 41375 34574 41384
rect 34808 41177 34836 42230
rect 34992 42090 35020 42638
rect 35084 42566 35112 42706
rect 35072 42560 35124 42566
rect 35072 42502 35124 42508
rect 35084 42401 35112 42502
rect 35070 42392 35126 42401
rect 35176 42362 35204 43114
rect 35070 42327 35072 42336
rect 35124 42327 35126 42336
rect 35164 42356 35216 42362
rect 35072 42298 35124 42304
rect 35164 42298 35216 42304
rect 34980 42084 35032 42090
rect 34980 42026 35032 42032
rect 34992 41682 35020 42026
rect 34980 41676 35032 41682
rect 34980 41618 35032 41624
rect 34888 41472 34940 41478
rect 34888 41414 34940 41420
rect 34794 41168 34850 41177
rect 34244 41132 34296 41138
rect 34794 41103 34850 41112
rect 34244 41074 34296 41080
rect 34900 41070 34928 41414
rect 34888 41064 34940 41070
rect 34888 41006 34940 41012
rect 34152 40996 34204 41002
rect 34152 40938 34204 40944
rect 33836 40548 33916 40576
rect 33784 40530 33836 40536
rect 33508 40520 33560 40526
rect 33508 40462 33560 40468
rect 33968 40520 34020 40526
rect 33968 40462 34020 40468
rect 34060 40520 34112 40526
rect 34060 40462 34112 40468
rect 33980 39642 34008 40462
rect 33968 39636 34020 39642
rect 33968 39578 34020 39584
rect 33692 39024 33744 39030
rect 33692 38966 33744 38972
rect 33704 37369 33732 38966
rect 33980 38962 34008 39578
rect 34072 39030 34100 40462
rect 34060 39024 34112 39030
rect 34060 38966 34112 38972
rect 33968 38956 34020 38962
rect 33968 38898 34020 38904
rect 34164 38826 34192 40938
rect 34612 40928 34664 40934
rect 34612 40870 34664 40876
rect 34624 40730 34652 40870
rect 34612 40724 34664 40730
rect 34612 40666 34664 40672
rect 34336 39500 34388 39506
rect 34336 39442 34388 39448
rect 34348 39302 34376 39442
rect 34612 39432 34664 39438
rect 34612 39374 34664 39380
rect 34336 39296 34388 39302
rect 34336 39238 34388 39244
rect 34624 39030 34652 39374
rect 34612 39024 34664 39030
rect 34612 38966 34664 38972
rect 33968 38820 34020 38826
rect 33968 38762 34020 38768
rect 34152 38820 34204 38826
rect 34152 38762 34204 38768
rect 33980 38486 34008 38762
rect 34336 38752 34388 38758
rect 34336 38694 34388 38700
rect 33968 38480 34020 38486
rect 33968 38422 34020 38428
rect 34244 38344 34296 38350
rect 34150 38312 34206 38321
rect 34244 38286 34296 38292
rect 34150 38247 34206 38256
rect 33784 37664 33836 37670
rect 33784 37606 33836 37612
rect 33690 37360 33746 37369
rect 33690 37295 33746 37304
rect 33796 37194 33824 37606
rect 33784 37188 33836 37194
rect 33784 37130 33836 37136
rect 33414 36000 33470 36009
rect 33414 35935 33470 35944
rect 31114 35864 31170 35873
rect 31114 35799 31170 35808
rect 33046 35864 33102 35873
rect 34164 35850 34192 38247
rect 34256 37942 34284 38286
rect 34348 38185 34376 38694
rect 34428 38548 34480 38554
rect 34428 38490 34480 38496
rect 34520 38548 34572 38554
rect 34520 38490 34572 38496
rect 34440 38321 34468 38490
rect 34426 38312 34482 38321
rect 34426 38247 34482 38256
rect 34334 38176 34390 38185
rect 34334 38111 34390 38120
rect 34244 37936 34296 37942
rect 34244 37878 34296 37884
rect 34336 37936 34388 37942
rect 34336 37878 34388 37884
rect 34348 37670 34376 37878
rect 34532 37670 34560 38490
rect 34704 38344 34756 38350
rect 34704 38286 34756 38292
rect 34336 37664 34388 37670
rect 34336 37606 34388 37612
rect 34520 37664 34572 37670
rect 34520 37606 34572 37612
rect 34518 37496 34574 37505
rect 34428 37460 34480 37466
rect 34518 37431 34520 37440
rect 34428 37402 34480 37408
rect 34572 37431 34574 37440
rect 34520 37402 34572 37408
rect 34440 37233 34468 37402
rect 34532 37330 34560 37402
rect 34520 37324 34572 37330
rect 34520 37266 34572 37272
rect 34716 37262 34744 38286
rect 34704 37256 34756 37262
rect 34426 37224 34482 37233
rect 34704 37198 34756 37204
rect 34426 37159 34482 37168
rect 34992 37126 35020 41618
rect 35256 41132 35308 41138
rect 35256 41074 35308 41080
rect 35072 40928 35124 40934
rect 35072 40870 35124 40876
rect 35084 40662 35112 40870
rect 35072 40656 35124 40662
rect 35072 40598 35124 40604
rect 35268 40118 35296 41074
rect 35256 40112 35308 40118
rect 35176 40072 35256 40100
rect 35072 39568 35124 39574
rect 35072 39510 35124 39516
rect 35084 39302 35112 39510
rect 35072 39296 35124 39302
rect 35072 39238 35124 39244
rect 35176 38350 35204 40072
rect 35256 40054 35308 40060
rect 35256 39840 35308 39846
rect 35256 39782 35308 39788
rect 35268 39545 35296 39782
rect 35254 39536 35310 39545
rect 35254 39471 35310 39480
rect 35164 38344 35216 38350
rect 35164 38286 35216 38292
rect 35256 38344 35308 38350
rect 35256 38286 35308 38292
rect 35176 37874 35204 38286
rect 35164 37868 35216 37874
rect 35164 37810 35216 37816
rect 35268 37466 35296 38286
rect 35360 37806 35388 45047
rect 40408 44736 40460 44742
rect 40408 44678 40460 44684
rect 36544 44532 36596 44538
rect 36544 44474 36596 44480
rect 35716 44396 35768 44402
rect 35716 44338 35768 44344
rect 35440 44328 35492 44334
rect 35440 44270 35492 44276
rect 35728 44282 35756 44338
rect 35452 43790 35480 44270
rect 35728 44254 35848 44282
rect 35532 44192 35584 44198
rect 35532 44134 35584 44140
rect 35440 43784 35492 43790
rect 35440 43726 35492 43732
rect 35452 42922 35480 43726
rect 35544 43722 35572 44134
rect 35532 43716 35584 43722
rect 35532 43658 35584 43664
rect 35452 42894 35572 42922
rect 35544 42838 35572 42894
rect 35532 42832 35584 42838
rect 35532 42774 35584 42780
rect 35716 42560 35768 42566
rect 35716 42502 35768 42508
rect 35728 42226 35756 42502
rect 35820 42226 35848 44254
rect 36556 43450 36584 44474
rect 38108 44464 38160 44470
rect 38292 44464 38344 44470
rect 38160 44412 38292 44418
rect 38108 44406 38344 44412
rect 39396 44464 39448 44470
rect 39396 44406 39448 44412
rect 37924 44396 37976 44402
rect 37924 44338 37976 44344
rect 38016 44396 38068 44402
rect 38120 44390 38332 44406
rect 38016 44338 38068 44344
rect 37740 44260 37792 44266
rect 37740 44202 37792 44208
rect 36636 44192 36688 44198
rect 36636 44134 36688 44140
rect 37464 44192 37516 44198
rect 37464 44134 37516 44140
rect 36648 43994 36676 44134
rect 36636 43988 36688 43994
rect 36636 43930 36688 43936
rect 37280 43988 37332 43994
rect 37280 43930 37332 43936
rect 36636 43852 36688 43858
rect 36636 43794 36688 43800
rect 36648 43654 36676 43794
rect 36636 43648 36688 43654
rect 36636 43590 36688 43596
rect 36648 43450 36676 43590
rect 36544 43444 36596 43450
rect 36544 43386 36596 43392
rect 36636 43444 36688 43450
rect 36636 43386 36688 43392
rect 36648 42770 36676 43386
rect 37096 43308 37148 43314
rect 37096 43250 37148 43256
rect 36818 43072 36874 43081
rect 36818 43007 36874 43016
rect 36832 42770 36860 43007
rect 36636 42764 36688 42770
rect 36636 42706 36688 42712
rect 36820 42764 36872 42770
rect 36820 42706 36872 42712
rect 35900 42560 35952 42566
rect 35900 42502 35952 42508
rect 35716 42220 35768 42226
rect 35716 42162 35768 42168
rect 35808 42220 35860 42226
rect 35808 42162 35860 42168
rect 35820 41414 35848 42162
rect 35912 42158 35940 42502
rect 36832 42362 36860 42706
rect 36820 42356 36872 42362
rect 36820 42298 36872 42304
rect 35900 42152 35952 42158
rect 35900 42094 35952 42100
rect 36268 42152 36320 42158
rect 36268 42094 36320 42100
rect 35900 41472 35952 41478
rect 35900 41414 35952 41420
rect 35728 41386 35848 41414
rect 35728 41138 35756 41386
rect 35808 41268 35860 41274
rect 35808 41210 35860 41216
rect 35716 41132 35768 41138
rect 35716 41074 35768 41080
rect 35440 40928 35492 40934
rect 35440 40870 35492 40876
rect 35452 39642 35480 40870
rect 35532 40656 35584 40662
rect 35532 40598 35584 40604
rect 35544 39914 35572 40598
rect 35820 40225 35848 41210
rect 35912 41138 35940 41414
rect 35900 41132 35952 41138
rect 35900 41074 35952 41080
rect 36280 41002 36308 42094
rect 37108 41750 37136 43250
rect 37292 42770 37320 43930
rect 37476 43314 37504 44134
rect 37556 43784 37608 43790
rect 37556 43726 37608 43732
rect 37464 43308 37516 43314
rect 37464 43250 37516 43256
rect 37280 42764 37332 42770
rect 37280 42706 37332 42712
rect 37568 42702 37596 43726
rect 37556 42696 37608 42702
rect 37556 42638 37608 42644
rect 37752 42634 37780 44202
rect 37936 43450 37964 44338
rect 37924 43444 37976 43450
rect 37924 43386 37976 43392
rect 38028 42702 38056 44338
rect 38292 44328 38344 44334
rect 38292 44270 38344 44276
rect 38108 44260 38160 44266
rect 38108 44202 38160 44208
rect 38120 43926 38148 44202
rect 38304 43994 38332 44270
rect 38752 44260 38804 44266
rect 38752 44202 38804 44208
rect 38292 43988 38344 43994
rect 38292 43930 38344 43936
rect 38108 43920 38160 43926
rect 38108 43862 38160 43868
rect 38660 43920 38712 43926
rect 38660 43862 38712 43868
rect 38672 42906 38700 43862
rect 38764 43178 38792 44202
rect 38844 44192 38896 44198
rect 38844 44134 38896 44140
rect 39028 44192 39080 44198
rect 39028 44134 39080 44140
rect 38856 43994 38884 44134
rect 38844 43988 38896 43994
rect 38844 43930 38896 43936
rect 38936 43852 38988 43858
rect 38936 43794 38988 43800
rect 38948 43314 38976 43794
rect 38936 43308 38988 43314
rect 38936 43250 38988 43256
rect 38752 43172 38804 43178
rect 38752 43114 38804 43120
rect 38568 42900 38620 42906
rect 38568 42842 38620 42848
rect 38660 42900 38712 42906
rect 38660 42842 38712 42848
rect 38016 42696 38068 42702
rect 38016 42638 38068 42644
rect 38384 42696 38436 42702
rect 38384 42638 38436 42644
rect 37740 42628 37792 42634
rect 37740 42570 37792 42576
rect 37832 42560 37884 42566
rect 37832 42502 37884 42508
rect 37844 42226 37872 42502
rect 37832 42220 37884 42226
rect 37832 42162 37884 42168
rect 37004 41744 37056 41750
rect 37004 41686 37056 41692
rect 37096 41744 37148 41750
rect 37096 41686 37148 41692
rect 36544 41608 36596 41614
rect 36544 41550 36596 41556
rect 36634 41576 36690 41585
rect 35900 40996 35952 41002
rect 35900 40938 35952 40944
rect 36268 40996 36320 41002
rect 36268 40938 36320 40944
rect 35912 40730 35940 40938
rect 35900 40724 35952 40730
rect 35900 40666 35952 40672
rect 36084 40520 36136 40526
rect 36084 40462 36136 40468
rect 35806 40216 35862 40225
rect 36096 40186 36124 40462
rect 36280 40186 36308 40938
rect 36450 40896 36506 40905
rect 36450 40831 36506 40840
rect 35806 40151 35862 40160
rect 36084 40180 36136 40186
rect 36084 40122 36136 40128
rect 36268 40180 36320 40186
rect 36268 40122 36320 40128
rect 36464 40050 36492 40831
rect 36556 40730 36584 41550
rect 36634 41511 36690 41520
rect 36544 40724 36596 40730
rect 36544 40666 36596 40672
rect 36452 40044 36504 40050
rect 36452 39986 36504 39992
rect 35532 39908 35584 39914
rect 35532 39850 35584 39856
rect 35992 39840 36044 39846
rect 35992 39782 36044 39788
rect 35440 39636 35492 39642
rect 35440 39578 35492 39584
rect 36004 39506 36032 39782
rect 36556 39574 36584 40666
rect 36544 39568 36596 39574
rect 36544 39510 36596 39516
rect 35992 39500 36044 39506
rect 35992 39442 36044 39448
rect 35808 39432 35860 39438
rect 35808 39374 35860 39380
rect 35440 39296 35492 39302
rect 35440 39238 35492 39244
rect 35452 38554 35480 39238
rect 35624 38820 35676 38826
rect 35624 38762 35676 38768
rect 35636 38554 35664 38762
rect 35440 38548 35492 38554
rect 35440 38490 35492 38496
rect 35624 38548 35676 38554
rect 35624 38490 35676 38496
rect 35348 37800 35400 37806
rect 35348 37742 35400 37748
rect 35440 37664 35492 37670
rect 35440 37606 35492 37612
rect 35452 37466 35480 37606
rect 35820 37466 35848 39374
rect 36648 37466 36676 41511
rect 37016 41177 37044 41686
rect 37108 41414 37136 41686
rect 38396 41682 38424 42638
rect 38580 41750 38608 42842
rect 38764 42090 38792 43114
rect 39040 42906 39068 44134
rect 39408 43858 39436 44406
rect 40420 44334 40448 44678
rect 50998 44636 51306 44645
rect 50998 44634 51004 44636
rect 51060 44634 51084 44636
rect 51140 44634 51164 44636
rect 51220 44634 51244 44636
rect 51300 44634 51306 44636
rect 51060 44582 51062 44634
rect 51242 44582 51244 44634
rect 50998 44580 51004 44582
rect 51060 44580 51084 44582
rect 51140 44580 51164 44582
rect 51220 44580 51244 44582
rect 51300 44580 51306 44582
rect 50998 44571 51306 44580
rect 41604 44532 41656 44538
rect 41604 44474 41656 44480
rect 42524 44532 42576 44538
rect 42524 44474 42576 44480
rect 39856 44328 39908 44334
rect 40408 44328 40460 44334
rect 39908 44288 39988 44316
rect 39856 44270 39908 44276
rect 39580 44192 39632 44198
rect 39580 44134 39632 44140
rect 39396 43852 39448 43858
rect 39396 43794 39448 43800
rect 39592 43722 39620 44134
rect 39960 43858 39988 44288
rect 40408 44270 40460 44276
rect 40500 44260 40552 44266
rect 40500 44202 40552 44208
rect 40868 44260 40920 44266
rect 40868 44202 40920 44208
rect 39948 43852 40000 43858
rect 39948 43794 40000 43800
rect 39580 43716 39632 43722
rect 39580 43658 39632 43664
rect 39304 43648 39356 43654
rect 39304 43590 39356 43596
rect 39316 42906 39344 43590
rect 39764 43240 39816 43246
rect 39764 43182 39816 43188
rect 39028 42900 39080 42906
rect 39028 42842 39080 42848
rect 39304 42900 39356 42906
rect 39304 42842 39356 42848
rect 39120 42764 39172 42770
rect 39120 42706 39172 42712
rect 38936 42356 38988 42362
rect 38936 42298 38988 42304
rect 38752 42084 38804 42090
rect 38752 42026 38804 42032
rect 38568 41744 38620 41750
rect 38568 41686 38620 41692
rect 38384 41676 38436 41682
rect 38384 41618 38436 41624
rect 37832 41608 37884 41614
rect 37832 41550 37884 41556
rect 37556 41472 37608 41478
rect 37556 41414 37608 41420
rect 37108 41386 37228 41414
rect 37094 41304 37150 41313
rect 37094 41239 37096 41248
rect 37148 41239 37150 41248
rect 37096 41210 37148 41216
rect 37002 41168 37058 41177
rect 37002 41103 37058 41112
rect 37200 41070 37228 41386
rect 37188 41064 37240 41070
rect 37094 41032 37150 41041
rect 37188 41006 37240 41012
rect 37094 40967 37096 40976
rect 37148 40967 37150 40976
rect 37096 40938 37148 40944
rect 36728 40180 36780 40186
rect 36728 40122 36780 40128
rect 36740 38418 36768 40122
rect 36820 39908 36872 39914
rect 36820 39850 36872 39856
rect 36832 39642 36860 39850
rect 36820 39636 36872 39642
rect 36820 39578 36872 39584
rect 36912 39636 36964 39642
rect 36912 39578 36964 39584
rect 36924 39522 36952 39578
rect 36832 39494 36952 39522
rect 36728 38412 36780 38418
rect 36728 38354 36780 38360
rect 35256 37460 35308 37466
rect 35256 37402 35308 37408
rect 35440 37460 35492 37466
rect 35440 37402 35492 37408
rect 35808 37460 35860 37466
rect 35808 37402 35860 37408
rect 36636 37460 36688 37466
rect 36636 37402 36688 37408
rect 35806 37360 35862 37369
rect 35806 37295 35862 37304
rect 34980 37120 35032 37126
rect 34980 37062 35032 37068
rect 35820 36854 35848 37295
rect 36084 37256 36136 37262
rect 36084 37198 36136 37204
rect 36096 37126 36124 37198
rect 36084 37120 36136 37126
rect 36176 37120 36228 37126
rect 36136 37080 36176 37108
rect 36084 37062 36136 37068
rect 36176 37062 36228 37068
rect 36832 36961 36860 39494
rect 36912 39432 36964 39438
rect 36912 39374 36964 39380
rect 36924 37330 36952 39374
rect 37004 38752 37056 38758
rect 37004 38694 37056 38700
rect 37016 38486 37044 38694
rect 37004 38480 37056 38486
rect 37004 38422 37056 38428
rect 37108 37874 37136 40938
rect 37200 40594 37228 41006
rect 37568 40662 37596 41414
rect 37844 41274 37872 41550
rect 37832 41268 37884 41274
rect 37832 41210 37884 41216
rect 37556 40656 37608 40662
rect 37556 40598 37608 40604
rect 37188 40588 37240 40594
rect 37188 40530 37240 40536
rect 37200 40050 37228 40530
rect 38396 40526 38424 41618
rect 38580 40730 38608 41686
rect 38948 41206 38976 42298
rect 39132 41274 39160 42706
rect 39304 42696 39356 42702
rect 39304 42638 39356 42644
rect 39316 42362 39344 42638
rect 39304 42356 39356 42362
rect 39304 42298 39356 42304
rect 39396 42084 39448 42090
rect 39396 42026 39448 42032
rect 39304 42016 39356 42022
rect 39304 41958 39356 41964
rect 39316 41818 39344 41958
rect 39304 41812 39356 41818
rect 39304 41754 39356 41760
rect 39120 41268 39172 41274
rect 39120 41210 39172 41216
rect 38936 41200 38988 41206
rect 38936 41142 38988 41148
rect 38568 40724 38620 40730
rect 38568 40666 38620 40672
rect 37648 40520 37700 40526
rect 37648 40462 37700 40468
rect 38384 40520 38436 40526
rect 38384 40462 38436 40468
rect 37278 40352 37334 40361
rect 37278 40287 37334 40296
rect 37188 40044 37240 40050
rect 37188 39986 37240 39992
rect 37200 38962 37228 39986
rect 37292 39846 37320 40287
rect 37370 40080 37426 40089
rect 37370 40015 37426 40024
rect 37280 39840 37332 39846
rect 37280 39782 37332 39788
rect 37384 39438 37412 40015
rect 37372 39432 37424 39438
rect 37372 39374 37424 39380
rect 37372 39296 37424 39302
rect 37372 39238 37424 39244
rect 37384 38962 37412 39238
rect 37188 38956 37240 38962
rect 37188 38898 37240 38904
rect 37372 38956 37424 38962
rect 37372 38898 37424 38904
rect 37200 37874 37228 38898
rect 37464 38752 37516 38758
rect 37464 38694 37516 38700
rect 37096 37868 37148 37874
rect 37096 37810 37148 37816
rect 37188 37868 37240 37874
rect 37188 37810 37240 37816
rect 37476 37738 37504 38694
rect 37464 37732 37516 37738
rect 37464 37674 37516 37680
rect 36912 37324 36964 37330
rect 36912 37266 36964 37272
rect 36818 36952 36874 36961
rect 36818 36887 36874 36896
rect 35808 36848 35860 36854
rect 35808 36790 35860 36796
rect 37660 36650 37688 40462
rect 38292 40044 38344 40050
rect 38292 39986 38344 39992
rect 38304 39506 38332 39986
rect 38292 39500 38344 39506
rect 38292 39442 38344 39448
rect 38304 38962 38332 39442
rect 38200 38956 38252 38962
rect 38200 38898 38252 38904
rect 38292 38956 38344 38962
rect 38292 38898 38344 38904
rect 38476 38956 38528 38962
rect 38476 38898 38528 38904
rect 38212 38758 38240 38898
rect 38016 38752 38068 38758
rect 38016 38694 38068 38700
rect 38200 38752 38252 38758
rect 38200 38694 38252 38700
rect 38028 38049 38056 38694
rect 38488 38554 38516 38898
rect 38476 38548 38528 38554
rect 38476 38490 38528 38496
rect 38014 38040 38070 38049
rect 38014 37975 38070 37984
rect 38580 37262 38608 40666
rect 39028 40656 39080 40662
rect 39028 40598 39080 40604
rect 38660 40384 38712 40390
rect 38660 40326 38712 40332
rect 38672 39817 38700 40326
rect 39040 39982 39068 40598
rect 39304 40520 39356 40526
rect 39304 40462 39356 40468
rect 39212 40384 39264 40390
rect 39212 40326 39264 40332
rect 39224 40186 39252 40326
rect 39212 40180 39264 40186
rect 39212 40122 39264 40128
rect 39028 39976 39080 39982
rect 39028 39918 39080 39924
rect 39040 39846 39068 39918
rect 39028 39840 39080 39846
rect 38658 39808 38714 39817
rect 39028 39782 39080 39788
rect 38658 39743 38714 39752
rect 38658 39264 38714 39273
rect 38658 39199 38714 39208
rect 38568 37256 38620 37262
rect 38568 37198 38620 37204
rect 38672 36854 38700 39199
rect 39316 39030 39344 40462
rect 39408 40186 39436 42026
rect 39488 41268 39540 41274
rect 39488 41210 39540 41216
rect 39396 40180 39448 40186
rect 39396 40122 39448 40128
rect 39408 39846 39436 40122
rect 39500 40050 39528 41210
rect 39776 41138 39804 43182
rect 39960 43110 39988 43794
rect 40224 43784 40276 43790
rect 40224 43726 40276 43732
rect 40132 43444 40184 43450
rect 40132 43386 40184 43392
rect 39948 43104 40000 43110
rect 39948 43046 40000 43052
rect 39960 42838 39988 43046
rect 39948 42832 40000 42838
rect 39948 42774 40000 42780
rect 39856 42016 39908 42022
rect 39856 41958 39908 41964
rect 39868 41614 39896 41958
rect 39856 41608 39908 41614
rect 39856 41550 39908 41556
rect 39764 41132 39816 41138
rect 39764 41074 39816 41080
rect 39856 40520 39908 40526
rect 39776 40468 39856 40474
rect 39776 40462 39908 40468
rect 39776 40446 39896 40462
rect 39488 40044 39540 40050
rect 39488 39986 39540 39992
rect 39396 39840 39448 39846
rect 39396 39782 39448 39788
rect 39672 39840 39724 39846
rect 39776 39828 39804 40446
rect 39724 39800 39804 39828
rect 39856 39840 39908 39846
rect 39672 39782 39724 39788
rect 39856 39782 39908 39788
rect 39408 39574 39436 39782
rect 39684 39642 39712 39782
rect 39672 39636 39724 39642
rect 39672 39578 39724 39584
rect 39396 39568 39448 39574
rect 39396 39510 39448 39516
rect 39120 39024 39172 39030
rect 39120 38966 39172 38972
rect 39304 39024 39356 39030
rect 39304 38966 39356 38972
rect 38936 38888 38988 38894
rect 38936 38830 38988 38836
rect 38752 38344 38804 38350
rect 38752 38286 38804 38292
rect 38764 37806 38792 38286
rect 38948 38049 38976 38830
rect 38934 38040 38990 38049
rect 38934 37975 38990 37984
rect 38948 37942 38976 37975
rect 38936 37936 38988 37942
rect 38936 37878 38988 37884
rect 38752 37800 38804 37806
rect 38752 37742 38804 37748
rect 38752 37460 38804 37466
rect 38752 37402 38804 37408
rect 38660 36848 38712 36854
rect 38660 36790 38712 36796
rect 38764 36786 38792 37402
rect 38948 37330 38976 37878
rect 39132 37466 39160 38966
rect 39684 38758 39712 39578
rect 39868 39574 39896 39782
rect 39856 39568 39908 39574
rect 39856 39510 39908 39516
rect 39672 38752 39724 38758
rect 39672 38694 39724 38700
rect 39856 38752 39908 38758
rect 39856 38694 39908 38700
rect 39868 38486 39896 38694
rect 39856 38480 39908 38486
rect 39856 38422 39908 38428
rect 39960 38468 39988 42774
rect 40040 42152 40092 42158
rect 40040 42094 40092 42100
rect 40052 40934 40080 42094
rect 40144 41206 40172 43386
rect 40236 41818 40264 43726
rect 40408 43172 40460 43178
rect 40408 43114 40460 43120
rect 40420 42906 40448 43114
rect 40408 42900 40460 42906
rect 40408 42842 40460 42848
rect 40512 42770 40540 44202
rect 40776 43784 40828 43790
rect 40776 43726 40828 43732
rect 40788 43314 40816 43726
rect 40776 43308 40828 43314
rect 40776 43250 40828 43256
rect 40880 43246 40908 44202
rect 41512 44192 41564 44198
rect 41512 44134 41564 44140
rect 41052 43988 41104 43994
rect 41052 43930 41104 43936
rect 40868 43240 40920 43246
rect 40868 43182 40920 43188
rect 40776 42900 40828 42906
rect 40776 42842 40828 42848
rect 40500 42764 40552 42770
rect 40500 42706 40552 42712
rect 40512 42566 40540 42706
rect 40500 42560 40552 42566
rect 40500 42502 40552 42508
rect 40316 42016 40368 42022
rect 40316 41958 40368 41964
rect 40224 41812 40276 41818
rect 40224 41754 40276 41760
rect 40132 41200 40184 41206
rect 40132 41142 40184 41148
rect 40040 40928 40092 40934
rect 40040 40870 40092 40876
rect 40052 40662 40080 40870
rect 40040 40656 40092 40662
rect 40040 40598 40092 40604
rect 40052 39642 40080 40598
rect 40132 40588 40184 40594
rect 40132 40530 40184 40536
rect 40144 40050 40172 40530
rect 40236 40050 40264 41754
rect 40328 40458 40356 41958
rect 40408 41608 40460 41614
rect 40408 41550 40460 41556
rect 40420 40934 40448 41550
rect 40684 41200 40736 41206
rect 40684 41142 40736 41148
rect 40408 40928 40460 40934
rect 40408 40870 40460 40876
rect 40696 40458 40724 41142
rect 40788 40662 40816 42842
rect 40880 42294 40908 43182
rect 41064 43110 41092 43930
rect 41420 43648 41472 43654
rect 41420 43590 41472 43596
rect 41328 43308 41380 43314
rect 41328 43250 41380 43256
rect 41052 43104 41104 43110
rect 41052 43046 41104 43052
rect 41064 42906 41092 43046
rect 41052 42900 41104 42906
rect 41052 42842 41104 42848
rect 41340 42770 41368 43250
rect 41432 42906 41460 43590
rect 41524 43178 41552 44134
rect 41512 43172 41564 43178
rect 41512 43114 41564 43120
rect 41420 42900 41472 42906
rect 41420 42842 41472 42848
rect 41328 42764 41380 42770
rect 41328 42706 41380 42712
rect 41616 42634 41644 44474
rect 42536 44402 42564 44474
rect 42524 44396 42576 44402
rect 42524 44338 42576 44344
rect 43076 44396 43128 44402
rect 43076 44338 43128 44344
rect 43996 44396 44048 44402
rect 43996 44338 44048 44344
rect 48228 44396 48280 44402
rect 48228 44338 48280 44344
rect 42248 44192 42300 44198
rect 42248 44134 42300 44140
rect 42340 44192 42392 44198
rect 42340 44134 42392 44140
rect 42432 44192 42484 44198
rect 42432 44134 42484 44140
rect 42260 43994 42288 44134
rect 42248 43988 42300 43994
rect 42248 43930 42300 43936
rect 41972 43784 42024 43790
rect 41972 43726 42024 43732
rect 41604 42628 41656 42634
rect 41604 42570 41656 42576
rect 40868 42288 40920 42294
rect 40868 42230 40920 42236
rect 41616 42226 41644 42570
rect 41604 42220 41656 42226
rect 41604 42162 41656 42168
rect 41696 42152 41748 42158
rect 41696 42094 41748 42100
rect 41708 41818 41736 42094
rect 41880 42084 41932 42090
rect 41880 42026 41932 42032
rect 41892 41993 41920 42026
rect 41878 41984 41934 41993
rect 41878 41919 41934 41928
rect 41696 41812 41748 41818
rect 41696 41754 41748 41760
rect 41328 41676 41380 41682
rect 41328 41618 41380 41624
rect 41340 41562 41368 41618
rect 41340 41534 41460 41562
rect 41432 41002 41460 41534
rect 41696 41472 41748 41478
rect 41696 41414 41748 41420
rect 41708 41002 41736 41414
rect 41984 41070 42012 43726
rect 42352 43450 42380 44134
rect 42444 43926 42472 44134
rect 42432 43920 42484 43926
rect 42432 43862 42484 43868
rect 42892 43920 42944 43926
rect 42892 43862 42944 43868
rect 42708 43784 42760 43790
rect 42708 43726 42760 43732
rect 42340 43444 42392 43450
rect 42340 43386 42392 43392
rect 42720 43382 42748 43726
rect 42708 43376 42760 43382
rect 42708 43318 42760 43324
rect 42616 43308 42668 43314
rect 42616 43250 42668 43256
rect 42064 42696 42116 42702
rect 42064 42638 42116 42644
rect 42076 42362 42104 42638
rect 42628 42566 42656 43250
rect 42524 42560 42576 42566
rect 42524 42502 42576 42508
rect 42616 42560 42668 42566
rect 42616 42502 42668 42508
rect 42064 42356 42116 42362
rect 42064 42298 42116 42304
rect 42432 42220 42484 42226
rect 42432 42162 42484 42168
rect 42444 41414 42472 42162
rect 42536 41818 42564 42502
rect 42628 42226 42656 42502
rect 42616 42220 42668 42226
rect 42616 42162 42668 42168
rect 42720 42158 42748 43318
rect 42904 43246 42932 43862
rect 43088 43450 43116 44338
rect 43812 44328 43864 44334
rect 43812 44270 43864 44276
rect 43824 43790 43852 44270
rect 43812 43784 43864 43790
rect 43812 43726 43864 43732
rect 43076 43444 43128 43450
rect 43076 43386 43128 43392
rect 43824 43382 43852 43726
rect 43812 43376 43864 43382
rect 43812 43318 43864 43324
rect 42892 43240 42944 43246
rect 42892 43182 42944 43188
rect 42904 42838 42932 43182
rect 43076 43104 43128 43110
rect 43076 43046 43128 43052
rect 43444 43104 43496 43110
rect 43444 43046 43496 43052
rect 42892 42832 42944 42838
rect 42892 42774 42944 42780
rect 42708 42152 42760 42158
rect 42708 42094 42760 42100
rect 43088 42022 43116 43046
rect 43456 42702 43484 43046
rect 43824 42906 43852 43318
rect 43904 43240 43956 43246
rect 43904 43182 43956 43188
rect 43812 42900 43864 42906
rect 43812 42842 43864 42848
rect 43720 42764 43772 42770
rect 43720 42706 43772 42712
rect 43444 42696 43496 42702
rect 43444 42638 43496 42644
rect 43352 42288 43404 42294
rect 43352 42230 43404 42236
rect 43076 42016 43128 42022
rect 43076 41958 43128 41964
rect 42524 41812 42576 41818
rect 42524 41754 42576 41760
rect 43364 41750 43392 42230
rect 43444 42084 43496 42090
rect 43444 42026 43496 42032
rect 43628 42084 43680 42090
rect 43628 42026 43680 42032
rect 43352 41744 43404 41750
rect 43352 41686 43404 41692
rect 42708 41608 42760 41614
rect 42708 41550 42760 41556
rect 42800 41608 42852 41614
rect 42800 41550 42852 41556
rect 43352 41608 43404 41614
rect 43352 41550 43404 41556
rect 42444 41386 42564 41414
rect 41972 41064 42024 41070
rect 41972 41006 42024 41012
rect 41420 40996 41472 41002
rect 41420 40938 41472 40944
rect 41604 40996 41656 41002
rect 41604 40938 41656 40944
rect 41696 40996 41748 41002
rect 41696 40938 41748 40944
rect 40960 40928 41012 40934
rect 40960 40870 41012 40876
rect 40776 40656 40828 40662
rect 40776 40598 40828 40604
rect 40972 40594 41000 40870
rect 41328 40656 41380 40662
rect 41328 40598 41380 40604
rect 40960 40588 41012 40594
rect 40960 40530 41012 40536
rect 40316 40452 40368 40458
rect 40316 40394 40368 40400
rect 40684 40452 40736 40458
rect 40684 40394 40736 40400
rect 40408 40384 40460 40390
rect 40408 40326 40460 40332
rect 40132 40044 40184 40050
rect 40132 39986 40184 39992
rect 40224 40044 40276 40050
rect 40224 39986 40276 39992
rect 40040 39636 40092 39642
rect 40040 39578 40092 39584
rect 40420 39506 40448 40326
rect 40408 39500 40460 39506
rect 40408 39442 40460 39448
rect 40224 39432 40276 39438
rect 40224 39374 40276 39380
rect 40132 39296 40184 39302
rect 40132 39238 40184 39244
rect 40144 39030 40172 39238
rect 40132 39024 40184 39030
rect 40132 38966 40184 38972
rect 40236 38962 40264 39374
rect 40224 38956 40276 38962
rect 40224 38898 40276 38904
rect 40040 38480 40092 38486
rect 39960 38440 40040 38468
rect 39960 38350 39988 38440
rect 40040 38422 40092 38428
rect 39948 38344 40000 38350
rect 39948 38286 40000 38292
rect 39960 37942 39988 38286
rect 39948 37936 40000 37942
rect 39948 37878 40000 37884
rect 40420 37874 40448 39442
rect 40696 39438 40724 40394
rect 40868 39976 40920 39982
rect 40868 39918 40920 39924
rect 40776 39636 40828 39642
rect 40776 39578 40828 39584
rect 40684 39432 40736 39438
rect 40684 39374 40736 39380
rect 40592 39296 40644 39302
rect 40592 39238 40644 39244
rect 40604 38962 40632 39238
rect 40592 38956 40644 38962
rect 40592 38898 40644 38904
rect 40788 38865 40816 39578
rect 40774 38856 40830 38865
rect 40774 38791 40830 38800
rect 40880 38554 40908 39918
rect 40972 39642 41000 40530
rect 40960 39636 41012 39642
rect 40960 39578 41012 39584
rect 41144 39500 41196 39506
rect 41144 39442 41196 39448
rect 41052 39296 41104 39302
rect 41052 39238 41104 39244
rect 41064 38894 41092 39238
rect 41052 38888 41104 38894
rect 41052 38830 41104 38836
rect 40868 38548 40920 38554
rect 40868 38490 40920 38496
rect 40868 38412 40920 38418
rect 40868 38354 40920 38360
rect 40776 38344 40828 38350
rect 40776 38286 40828 38292
rect 40788 38214 40816 38286
rect 40776 38208 40828 38214
rect 40776 38150 40828 38156
rect 40408 37868 40460 37874
rect 40408 37810 40460 37816
rect 39948 37664 40000 37670
rect 39948 37606 40000 37612
rect 39120 37460 39172 37466
rect 39120 37402 39172 37408
rect 39960 37330 39988 37606
rect 40788 37466 40816 38150
rect 40776 37460 40828 37466
rect 40776 37402 40828 37408
rect 38936 37324 38988 37330
rect 38936 37266 38988 37272
rect 39948 37324 40000 37330
rect 39948 37266 40000 37272
rect 40880 37262 40908 38354
rect 41156 37874 41184 39442
rect 41236 38956 41288 38962
rect 41236 38898 41288 38904
rect 41052 37868 41104 37874
rect 41052 37810 41104 37816
rect 41144 37868 41196 37874
rect 41144 37810 41196 37816
rect 40960 37732 41012 37738
rect 41064 37720 41092 37810
rect 41144 37732 41196 37738
rect 41064 37692 41144 37720
rect 40960 37674 41012 37680
rect 41144 37674 41196 37680
rect 40972 37466 41000 37674
rect 40960 37460 41012 37466
rect 40960 37402 41012 37408
rect 41248 37262 41276 38898
rect 41340 38418 41368 40598
rect 41616 40186 41644 40938
rect 41984 40594 42012 41006
rect 42248 40996 42300 41002
rect 42248 40938 42300 40944
rect 41972 40588 42024 40594
rect 41972 40530 42024 40536
rect 41604 40180 41656 40186
rect 41604 40122 41656 40128
rect 41880 40180 41932 40186
rect 41880 40122 41932 40128
rect 41892 39914 41920 40122
rect 41420 39908 41472 39914
rect 41420 39850 41472 39856
rect 41880 39908 41932 39914
rect 41880 39850 41932 39856
rect 41432 38554 41460 39850
rect 41604 39432 41656 39438
rect 41604 39374 41656 39380
rect 41512 38752 41564 38758
rect 41512 38694 41564 38700
rect 41420 38548 41472 38554
rect 41420 38490 41472 38496
rect 41328 38412 41380 38418
rect 41328 38354 41380 38360
rect 41340 38214 41368 38354
rect 41524 38282 41552 38694
rect 41616 38350 41644 39374
rect 41788 39296 41840 39302
rect 41788 39238 41840 39244
rect 41800 39098 41828 39238
rect 41788 39092 41840 39098
rect 41788 39034 41840 39040
rect 41892 38894 41920 39850
rect 42260 39642 42288 40938
rect 42432 39976 42484 39982
rect 42432 39918 42484 39924
rect 42248 39636 42300 39642
rect 42248 39578 42300 39584
rect 41880 38888 41932 38894
rect 41694 38856 41750 38865
rect 41880 38830 41932 38836
rect 41694 38791 41696 38800
rect 41748 38791 41750 38800
rect 41696 38762 41748 38768
rect 42260 38758 42288 39578
rect 42444 39302 42472 39918
rect 42432 39296 42484 39302
rect 42432 39238 42484 39244
rect 42248 38752 42300 38758
rect 42248 38694 42300 38700
rect 41604 38344 41656 38350
rect 41604 38286 41656 38292
rect 41512 38276 41564 38282
rect 41512 38218 41564 38224
rect 41328 38208 41380 38214
rect 41328 38150 41380 38156
rect 41328 37868 41380 37874
rect 41328 37810 41380 37816
rect 41340 37330 41368 37810
rect 42260 37806 42288 38694
rect 42536 38350 42564 41386
rect 42720 41206 42748 41550
rect 42708 41200 42760 41206
rect 42708 41142 42760 41148
rect 42812 41070 42840 41550
rect 43076 41132 43128 41138
rect 43076 41074 43128 41080
rect 42800 41064 42852 41070
rect 42800 41006 42852 41012
rect 43088 40934 43116 41074
rect 43168 40996 43220 41002
rect 43168 40938 43220 40944
rect 42800 40928 42852 40934
rect 42800 40870 42852 40876
rect 42892 40928 42944 40934
rect 42892 40870 42944 40876
rect 43076 40928 43128 40934
rect 43076 40870 43128 40876
rect 42616 39296 42668 39302
rect 42616 39238 42668 39244
rect 42628 38554 42656 39238
rect 42812 38944 42840 40870
rect 42904 39846 42932 40870
rect 43180 40746 43208 40938
rect 43088 40718 43208 40746
rect 43088 40050 43116 40718
rect 43364 40390 43392 41550
rect 43352 40384 43404 40390
rect 43352 40326 43404 40332
rect 43076 40044 43128 40050
rect 43076 39986 43128 39992
rect 42892 39840 42944 39846
rect 42892 39782 42944 39788
rect 43088 39642 43116 39986
rect 43260 39840 43312 39846
rect 43260 39782 43312 39788
rect 43076 39636 43128 39642
rect 43076 39578 43128 39584
rect 43088 39506 43116 39578
rect 43076 39500 43128 39506
rect 43076 39442 43128 39448
rect 42892 38956 42944 38962
rect 42812 38916 42892 38944
rect 42892 38898 42944 38904
rect 42616 38548 42668 38554
rect 42616 38490 42668 38496
rect 42708 38548 42760 38554
rect 42708 38490 42760 38496
rect 42524 38344 42576 38350
rect 42524 38286 42576 38292
rect 42720 37942 42748 38490
rect 43272 38418 43300 39782
rect 43364 38894 43392 40326
rect 43456 39574 43484 42026
rect 43640 41414 43668 42026
rect 43548 41386 43668 41414
rect 43548 39846 43576 41386
rect 43732 40526 43760 42706
rect 43916 42566 43944 43182
rect 43904 42560 43956 42566
rect 43904 42502 43956 42508
rect 43916 42294 43944 42502
rect 43904 42288 43956 42294
rect 43904 42230 43956 42236
rect 44008 42226 44036 44338
rect 47400 44328 47452 44334
rect 47400 44270 47452 44276
rect 44456 44192 44508 44198
rect 44456 44134 44508 44140
rect 45376 44192 45428 44198
rect 45376 44134 45428 44140
rect 46940 44192 46992 44198
rect 46940 44134 46992 44140
rect 44180 42696 44232 42702
rect 44180 42638 44232 42644
rect 44088 42560 44140 42566
rect 44088 42502 44140 42508
rect 43996 42220 44048 42226
rect 43996 42162 44048 42168
rect 43720 40520 43772 40526
rect 43720 40462 43772 40468
rect 43732 40050 43760 40462
rect 43720 40044 43772 40050
rect 43720 39986 43772 39992
rect 43536 39840 43588 39846
rect 43536 39782 43588 39788
rect 43444 39568 43496 39574
rect 43444 39510 43496 39516
rect 43812 39568 43864 39574
rect 43812 39510 43864 39516
rect 43824 39438 43852 39510
rect 43444 39432 43496 39438
rect 43444 39374 43496 39380
rect 43812 39432 43864 39438
rect 43812 39374 43864 39380
rect 43456 39098 43484 39374
rect 43444 39092 43496 39098
rect 43444 39034 43496 39040
rect 43628 39024 43680 39030
rect 43628 38966 43680 38972
rect 43352 38888 43404 38894
rect 43640 38865 43668 38966
rect 44008 38962 44036 42162
rect 44100 42158 44128 42502
rect 44192 42158 44220 42638
rect 44088 42152 44140 42158
rect 44088 42094 44140 42100
rect 44180 42152 44232 42158
rect 44180 42094 44232 42100
rect 44468 42022 44496 44134
rect 45388 43926 45416 44134
rect 45376 43920 45428 43926
rect 45376 43862 45428 43868
rect 46020 43920 46072 43926
rect 46020 43862 46072 43868
rect 45100 43784 45152 43790
rect 45100 43726 45152 43732
rect 44916 43104 44968 43110
rect 44916 43046 44968 43052
rect 44928 42906 44956 43046
rect 44916 42900 44968 42906
rect 44916 42842 44968 42848
rect 44456 42016 44508 42022
rect 44456 41958 44508 41964
rect 44824 42016 44876 42022
rect 44824 41958 44876 41964
rect 44836 41857 44864 41958
rect 44822 41848 44878 41857
rect 44822 41783 44878 41792
rect 45112 41682 45140 43726
rect 46032 43178 46060 43862
rect 46020 43172 46072 43178
rect 46020 43114 46072 43120
rect 46032 42906 46060 43114
rect 46952 42906 46980 44134
rect 47412 43994 47440 44270
rect 47400 43988 47452 43994
rect 47400 43930 47452 43936
rect 48044 43852 48096 43858
rect 48044 43794 48096 43800
rect 47216 43784 47268 43790
rect 47216 43726 47268 43732
rect 47584 43784 47636 43790
rect 47584 43726 47636 43732
rect 47228 43314 47256 43726
rect 47308 43648 47360 43654
rect 47308 43590 47360 43596
rect 47320 43314 47348 43590
rect 47216 43308 47268 43314
rect 47216 43250 47268 43256
rect 47308 43308 47360 43314
rect 47308 43250 47360 43256
rect 47228 42906 47256 43250
rect 47400 43172 47452 43178
rect 47400 43114 47452 43120
rect 46020 42900 46072 42906
rect 46020 42842 46072 42848
rect 46940 42900 46992 42906
rect 46940 42842 46992 42848
rect 47216 42900 47268 42906
rect 47216 42842 47268 42848
rect 45652 42696 45704 42702
rect 45652 42638 45704 42644
rect 45468 42220 45520 42226
rect 45468 42162 45520 42168
rect 45480 41750 45508 42162
rect 45558 42120 45614 42129
rect 45558 42055 45614 42064
rect 45572 42022 45600 42055
rect 45560 42016 45612 42022
rect 45560 41958 45612 41964
rect 45468 41744 45520 41750
rect 45468 41686 45520 41692
rect 45100 41676 45152 41682
rect 45100 41618 45152 41624
rect 44456 41608 44508 41614
rect 44456 41550 44508 41556
rect 44468 40644 44496 41550
rect 45008 41064 45060 41070
rect 45008 41006 45060 41012
rect 44732 40656 44784 40662
rect 44468 40616 44732 40644
rect 44732 40598 44784 40604
rect 44088 40044 44140 40050
rect 44088 39986 44140 39992
rect 43996 38956 44048 38962
rect 43996 38898 44048 38904
rect 43352 38830 43404 38836
rect 43626 38856 43682 38865
rect 43626 38791 43682 38800
rect 43260 38412 43312 38418
rect 43260 38354 43312 38360
rect 44100 38298 44128 39986
rect 44548 39432 44600 39438
rect 44548 39374 44600 39380
rect 44560 38865 44588 39374
rect 44824 39296 44876 39302
rect 44824 39238 44876 39244
rect 44546 38856 44602 38865
rect 44546 38791 44602 38800
rect 44180 38752 44232 38758
rect 44180 38694 44232 38700
rect 44008 38282 44128 38298
rect 43996 38276 44128 38282
rect 44048 38270 44128 38276
rect 43996 38218 44048 38224
rect 43812 38208 43864 38214
rect 43812 38150 43864 38156
rect 42708 37936 42760 37942
rect 42708 37878 42760 37884
rect 42248 37800 42300 37806
rect 42248 37742 42300 37748
rect 43824 37670 43852 38150
rect 44100 37874 44128 38270
rect 44192 38010 44220 38694
rect 44560 38486 44588 38791
rect 44548 38480 44600 38486
rect 44548 38422 44600 38428
rect 44456 38344 44508 38350
rect 44456 38286 44508 38292
rect 44468 38010 44496 38286
rect 44180 38004 44232 38010
rect 44180 37946 44232 37952
rect 44456 38004 44508 38010
rect 44456 37946 44508 37952
rect 44088 37868 44140 37874
rect 44088 37810 44140 37816
rect 44560 37738 44588 38422
rect 44836 38214 44864 39238
rect 44824 38208 44876 38214
rect 44824 38150 44876 38156
rect 44836 37806 44864 38150
rect 45020 37874 45048 41006
rect 45112 41002 45140 41618
rect 45664 41154 45692 42638
rect 46032 42090 46060 42842
rect 46572 42764 46624 42770
rect 46572 42706 46624 42712
rect 46388 42696 46440 42702
rect 46388 42638 46440 42644
rect 46020 42084 46072 42090
rect 46020 42026 46072 42032
rect 46032 41750 46060 42026
rect 46400 41818 46428 42638
rect 46388 41812 46440 41818
rect 46388 41754 46440 41760
rect 46020 41744 46072 41750
rect 46020 41686 46072 41692
rect 46032 41414 46060 41686
rect 46032 41386 46244 41414
rect 46112 41200 46164 41206
rect 45664 41126 45784 41154
rect 46112 41142 46164 41148
rect 45100 40996 45152 41002
rect 45100 40938 45152 40944
rect 45468 40996 45520 41002
rect 45468 40938 45520 40944
rect 45480 40594 45508 40938
rect 45756 40662 45784 41126
rect 46124 40934 46152 41142
rect 46112 40928 46164 40934
rect 46112 40870 46164 40876
rect 45744 40656 45796 40662
rect 45744 40598 45796 40604
rect 46216 40594 46244 41386
rect 46296 40928 46348 40934
rect 46296 40870 46348 40876
rect 45468 40588 45520 40594
rect 45468 40530 45520 40536
rect 46204 40588 46256 40594
rect 46204 40530 46256 40536
rect 45376 39976 45428 39982
rect 45376 39918 45428 39924
rect 45192 39840 45244 39846
rect 45192 39782 45244 39788
rect 45204 39681 45232 39782
rect 45190 39672 45246 39681
rect 45388 39642 45416 39918
rect 46216 39914 46244 40530
rect 46308 40186 46336 40870
rect 46400 40662 46428 41754
rect 46480 40996 46532 41002
rect 46480 40938 46532 40944
rect 46388 40656 46440 40662
rect 46388 40598 46440 40604
rect 46296 40180 46348 40186
rect 46296 40122 46348 40128
rect 46204 39908 46256 39914
rect 46204 39850 46256 39856
rect 45466 39672 45522 39681
rect 45190 39607 45246 39616
rect 45376 39636 45428 39642
rect 45466 39607 45522 39616
rect 45376 39578 45428 39584
rect 45284 38888 45336 38894
rect 45284 38830 45336 38836
rect 45192 38820 45244 38826
rect 45192 38762 45244 38768
rect 45204 38554 45232 38762
rect 45192 38548 45244 38554
rect 45192 38490 45244 38496
rect 45296 38418 45324 38830
rect 45480 38826 45508 39607
rect 46216 39574 46244 39850
rect 46492 39846 46520 40938
rect 46480 39840 46532 39846
rect 46480 39782 46532 39788
rect 46204 39568 46256 39574
rect 46204 39510 46256 39516
rect 45560 38956 45612 38962
rect 45560 38898 45612 38904
rect 45468 38820 45520 38826
rect 45468 38762 45520 38768
rect 45572 38758 45600 38898
rect 46584 38842 46612 42706
rect 46940 42220 46992 42226
rect 46940 42162 46992 42168
rect 46952 42022 46980 42162
rect 47032 42084 47084 42090
rect 47032 42026 47084 42032
rect 46848 42016 46900 42022
rect 46848 41958 46900 41964
rect 46940 42016 46992 42022
rect 46940 41958 46992 41964
rect 46860 41750 46888 41958
rect 47044 41818 47072 42026
rect 47228 41818 47256 42842
rect 47412 42226 47440 43114
rect 47492 42696 47544 42702
rect 47492 42638 47544 42644
rect 47400 42220 47452 42226
rect 47400 42162 47452 42168
rect 47032 41812 47084 41818
rect 47032 41754 47084 41760
rect 47216 41812 47268 41818
rect 47216 41754 47268 41760
rect 46848 41744 46900 41750
rect 46848 41686 46900 41692
rect 46664 40928 46716 40934
rect 46664 40870 46716 40876
rect 46676 39914 46704 40870
rect 47412 40458 47440 42162
rect 47504 41750 47532 42638
rect 47596 42634 47624 43726
rect 47768 43648 47820 43654
rect 47768 43590 47820 43596
rect 47780 42702 47808 43590
rect 47768 42696 47820 42702
rect 47768 42638 47820 42644
rect 47584 42628 47636 42634
rect 47584 42570 47636 42576
rect 47492 41744 47544 41750
rect 47492 41686 47544 41692
rect 47504 41002 47532 41686
rect 47596 41614 47624 42570
rect 47676 42560 47728 42566
rect 47676 42502 47728 42508
rect 47688 42226 47716 42502
rect 47676 42220 47728 42226
rect 47676 42162 47728 42168
rect 47584 41608 47636 41614
rect 47584 41550 47636 41556
rect 47780 41478 47808 42638
rect 47860 41744 47912 41750
rect 47860 41686 47912 41692
rect 47768 41472 47820 41478
rect 47768 41414 47820 41420
rect 47780 41120 47808 41414
rect 47872 41274 47900 41686
rect 47952 41676 48004 41682
rect 47952 41618 48004 41624
rect 47860 41268 47912 41274
rect 47860 41210 47912 41216
rect 47964 41138 47992 41618
rect 47860 41132 47912 41138
rect 47780 41092 47860 41120
rect 47860 41074 47912 41080
rect 47952 41132 48004 41138
rect 47952 41074 48004 41080
rect 47492 40996 47544 41002
rect 47492 40938 47544 40944
rect 47676 40588 47728 40594
rect 47676 40530 47728 40536
rect 47768 40588 47820 40594
rect 47768 40530 47820 40536
rect 47400 40452 47452 40458
rect 47400 40394 47452 40400
rect 47412 40050 47440 40394
rect 47400 40044 47452 40050
rect 47400 39986 47452 39992
rect 46664 39908 46716 39914
rect 46664 39850 46716 39856
rect 46676 39642 46704 39850
rect 47400 39840 47452 39846
rect 47400 39782 47452 39788
rect 47412 39642 47440 39782
rect 46664 39636 46716 39642
rect 46664 39578 46716 39584
rect 47400 39636 47452 39642
rect 47400 39578 47452 39584
rect 47492 39432 47544 39438
rect 47492 39374 47544 39380
rect 47504 39098 47532 39374
rect 47688 39098 47716 40530
rect 47780 40390 47808 40530
rect 47872 40526 47900 41074
rect 48056 41002 48084 43794
rect 48136 43172 48188 43178
rect 48136 43114 48188 43120
rect 48148 42770 48176 43114
rect 48240 42770 48268 44338
rect 50344 44260 50396 44266
rect 50344 44202 50396 44208
rect 48688 43784 48740 43790
rect 48688 43726 48740 43732
rect 48700 43314 48728 43726
rect 49424 43648 49476 43654
rect 49424 43590 49476 43596
rect 48688 43308 48740 43314
rect 48688 43250 48740 43256
rect 48700 42906 48728 43250
rect 49148 43172 49200 43178
rect 49148 43114 49200 43120
rect 49160 42906 49188 43114
rect 49436 42906 49464 43590
rect 49976 43240 50028 43246
rect 49976 43182 50028 43188
rect 48688 42900 48740 42906
rect 48688 42842 48740 42848
rect 49148 42900 49200 42906
rect 49148 42842 49200 42848
rect 49424 42900 49476 42906
rect 49424 42842 49476 42848
rect 49988 42770 50016 43182
rect 48136 42764 48188 42770
rect 48136 42706 48188 42712
rect 48228 42764 48280 42770
rect 48228 42706 48280 42712
rect 49976 42764 50028 42770
rect 49976 42706 50028 42712
rect 48148 42090 48176 42706
rect 48136 42084 48188 42090
rect 48136 42026 48188 42032
rect 48240 41546 48268 42706
rect 48688 42696 48740 42702
rect 48688 42638 48740 42644
rect 49516 42696 49568 42702
rect 49516 42638 49568 42644
rect 48700 42226 48728 42638
rect 48780 42560 48832 42566
rect 48780 42502 48832 42508
rect 48688 42220 48740 42226
rect 48688 42162 48740 42168
rect 48596 41676 48648 41682
rect 48596 41618 48648 41624
rect 48228 41540 48280 41546
rect 48228 41482 48280 41488
rect 48044 40996 48096 41002
rect 48044 40938 48096 40944
rect 47860 40520 47912 40526
rect 47860 40462 47912 40468
rect 47768 40384 47820 40390
rect 47768 40326 47820 40332
rect 47780 40118 47808 40326
rect 47768 40112 47820 40118
rect 47768 40054 47820 40060
rect 47780 39438 47808 40054
rect 47768 39432 47820 39438
rect 47768 39374 47820 39380
rect 47492 39092 47544 39098
rect 47492 39034 47544 39040
rect 47676 39092 47728 39098
rect 47676 39034 47728 39040
rect 46662 38856 46718 38865
rect 46204 38820 46256 38826
rect 46584 38814 46662 38842
rect 46662 38791 46664 38800
rect 46204 38762 46256 38768
rect 46716 38791 46718 38800
rect 47490 38856 47546 38865
rect 47780 38842 47808 39374
rect 47490 38791 47492 38800
rect 46664 38762 46716 38768
rect 47544 38791 47546 38800
rect 47688 38814 47808 38842
rect 47492 38762 47544 38768
rect 45376 38752 45428 38758
rect 45376 38694 45428 38700
rect 45560 38752 45612 38758
rect 45560 38694 45612 38700
rect 45284 38412 45336 38418
rect 45284 38354 45336 38360
rect 45008 37868 45060 37874
rect 45008 37810 45060 37816
rect 44824 37800 44876 37806
rect 44824 37742 44876 37748
rect 44548 37732 44600 37738
rect 44548 37674 44600 37680
rect 45388 37670 45416 38694
rect 46216 38554 46244 38762
rect 47124 38752 47176 38758
rect 47124 38694 47176 38700
rect 46204 38548 46256 38554
rect 46204 38490 46256 38496
rect 46572 38344 46624 38350
rect 46572 38286 46624 38292
rect 46756 38344 46808 38350
rect 46756 38286 46808 38292
rect 42064 37664 42116 37670
rect 43812 37664 43864 37670
rect 42064 37606 42116 37612
rect 43810 37632 43812 37641
rect 45376 37664 45428 37670
rect 43864 37632 43866 37641
rect 42076 37330 42104 37606
rect 45376 37606 45428 37612
rect 43810 37567 43866 37576
rect 46584 37466 46612 38286
rect 46768 38010 46796 38286
rect 46756 38004 46808 38010
rect 46756 37946 46808 37952
rect 46572 37460 46624 37466
rect 46572 37402 46624 37408
rect 46768 37398 46796 37946
rect 47136 37874 47164 38694
rect 47688 38418 47716 38814
rect 47768 38752 47820 38758
rect 47768 38694 47820 38700
rect 47780 38554 47808 38694
rect 47768 38548 47820 38554
rect 47768 38490 47820 38496
rect 47308 38412 47360 38418
rect 47308 38354 47360 38360
rect 47676 38412 47728 38418
rect 47676 38354 47728 38360
rect 47124 37868 47176 37874
rect 47124 37810 47176 37816
rect 46756 37392 46808 37398
rect 46756 37334 46808 37340
rect 41328 37324 41380 37330
rect 41328 37266 41380 37272
rect 42064 37324 42116 37330
rect 42064 37266 42116 37272
rect 47136 37262 47164 37810
rect 47320 37262 47348 38354
rect 47492 38208 47544 38214
rect 47492 38150 47544 38156
rect 47504 37466 47532 38150
rect 47872 37874 47900 40462
rect 48056 40186 48084 40938
rect 48240 40594 48268 41482
rect 48608 41274 48636 41618
rect 48596 41268 48648 41274
rect 48596 41210 48648 41216
rect 48792 41138 48820 42502
rect 49056 42220 49108 42226
rect 49056 42162 49108 42168
rect 49068 41818 49096 42162
rect 49528 41818 49556 42638
rect 49056 41812 49108 41818
rect 49056 41754 49108 41760
rect 49516 41812 49568 41818
rect 49516 41754 49568 41760
rect 48780 41132 48832 41138
rect 48780 41074 48832 41080
rect 49068 40769 49096 41754
rect 49988 41546 50016 42706
rect 50356 42702 50384 44202
rect 51918 44092 52226 44101
rect 51918 44090 51924 44092
rect 51980 44090 52004 44092
rect 52060 44090 52084 44092
rect 52140 44090 52164 44092
rect 52220 44090 52226 44092
rect 51980 44038 51982 44090
rect 52162 44038 52164 44090
rect 51918 44036 51924 44038
rect 51980 44036 52004 44038
rect 52060 44036 52084 44038
rect 52140 44036 52164 44038
rect 52220 44036 52226 44038
rect 51918 44027 52226 44036
rect 50998 43548 51306 43557
rect 50998 43546 51004 43548
rect 51060 43546 51084 43548
rect 51140 43546 51164 43548
rect 51220 43546 51244 43548
rect 51300 43546 51306 43548
rect 51060 43494 51062 43546
rect 51242 43494 51244 43546
rect 50998 43492 51004 43494
rect 51060 43492 51084 43494
rect 51140 43492 51164 43494
rect 51220 43492 51244 43494
rect 51300 43492 51306 43494
rect 50998 43483 51306 43492
rect 51724 43240 51776 43246
rect 51724 43182 51776 43188
rect 51540 43104 51592 43110
rect 51540 43046 51592 43052
rect 50252 42696 50304 42702
rect 50252 42638 50304 42644
rect 50344 42696 50396 42702
rect 50344 42638 50396 42644
rect 50804 42696 50856 42702
rect 50804 42638 50856 42644
rect 50264 41818 50292 42638
rect 50620 42084 50672 42090
rect 50620 42026 50672 42032
rect 50252 41812 50304 41818
rect 50252 41754 50304 41760
rect 49976 41540 50028 41546
rect 49976 41482 50028 41488
rect 50632 41138 50660 42026
rect 50816 41614 50844 42638
rect 50998 42460 51306 42469
rect 50998 42458 51004 42460
rect 51060 42458 51084 42460
rect 51140 42458 51164 42460
rect 51220 42458 51244 42460
rect 51300 42458 51306 42460
rect 51060 42406 51062 42458
rect 51242 42406 51244 42458
rect 50998 42404 51004 42406
rect 51060 42404 51084 42406
rect 51140 42404 51164 42406
rect 51220 42404 51244 42406
rect 51300 42404 51306 42406
rect 50998 42395 51306 42404
rect 51356 42220 51408 42226
rect 51356 42162 51408 42168
rect 51368 41682 51396 42162
rect 51552 41818 51580 43046
rect 51632 42764 51684 42770
rect 51632 42706 51684 42712
rect 51644 42362 51672 42706
rect 51736 42566 51764 43182
rect 52368 43172 52420 43178
rect 52368 43114 52420 43120
rect 51816 43104 51868 43110
rect 51816 43046 51868 43052
rect 51828 42838 51856 43046
rect 51918 43004 52226 43013
rect 51918 43002 51924 43004
rect 51980 43002 52004 43004
rect 52060 43002 52084 43004
rect 52140 43002 52164 43004
rect 52220 43002 52226 43004
rect 51980 42950 51982 43002
rect 52162 42950 52164 43002
rect 51918 42948 51924 42950
rect 51980 42948 52004 42950
rect 52060 42948 52084 42950
rect 52140 42948 52164 42950
rect 52220 42948 52226 42950
rect 51918 42939 52226 42948
rect 51816 42832 51868 42838
rect 51816 42774 51868 42780
rect 51724 42560 51776 42566
rect 51724 42502 51776 42508
rect 51736 42362 51764 42502
rect 51632 42356 51684 42362
rect 51632 42298 51684 42304
rect 51724 42356 51776 42362
rect 51724 42298 51776 42304
rect 51828 42090 51856 42774
rect 52380 42634 52408 43114
rect 60004 42764 60056 42770
rect 60004 42706 60056 42712
rect 54024 42696 54076 42702
rect 54024 42638 54076 42644
rect 54116 42696 54168 42702
rect 54116 42638 54168 42644
rect 52368 42628 52420 42634
rect 52368 42570 52420 42576
rect 53104 42560 53156 42566
rect 53104 42502 53156 42508
rect 53116 42158 53144 42502
rect 54036 42158 54064 42638
rect 53104 42152 53156 42158
rect 53104 42094 53156 42100
rect 54024 42152 54076 42158
rect 54024 42094 54076 42100
rect 51816 42084 51868 42090
rect 51816 42026 51868 42032
rect 51828 41818 51856 42026
rect 52276 42016 52328 42022
rect 52276 41958 52328 41964
rect 52460 42016 52512 42022
rect 52460 41958 52512 41964
rect 53196 42016 53248 42022
rect 53196 41958 53248 41964
rect 54024 42016 54076 42022
rect 54024 41958 54076 41964
rect 51918 41916 52226 41925
rect 51918 41914 51924 41916
rect 51980 41914 52004 41916
rect 52060 41914 52084 41916
rect 52140 41914 52164 41916
rect 52220 41914 52226 41916
rect 51980 41862 51982 41914
rect 52162 41862 52164 41914
rect 51918 41860 51924 41862
rect 51980 41860 52004 41862
rect 52060 41860 52084 41862
rect 52140 41860 52164 41862
rect 52220 41860 52226 41862
rect 51918 41851 52226 41860
rect 51540 41812 51592 41818
rect 51540 41754 51592 41760
rect 51816 41812 51868 41818
rect 51816 41754 51868 41760
rect 51448 41744 51500 41750
rect 51448 41686 51500 41692
rect 51356 41676 51408 41682
rect 51356 41618 51408 41624
rect 50804 41608 50856 41614
rect 50804 41550 50856 41556
rect 50896 41540 50948 41546
rect 50896 41482 50948 41488
rect 49332 41132 49384 41138
rect 49332 41074 49384 41080
rect 50620 41132 50672 41138
rect 50620 41074 50672 41080
rect 49054 40760 49110 40769
rect 49110 40718 49188 40746
rect 49054 40695 49110 40704
rect 48228 40588 48280 40594
rect 48228 40530 48280 40536
rect 48504 40520 48556 40526
rect 48504 40462 48556 40468
rect 48228 40452 48280 40458
rect 48228 40394 48280 40400
rect 48044 40180 48096 40186
rect 48044 40122 48096 40128
rect 48240 38418 48268 40394
rect 48516 40186 48544 40462
rect 49056 40384 49108 40390
rect 49056 40326 49108 40332
rect 48504 40180 48556 40186
rect 48504 40122 48556 40128
rect 49068 39982 49096 40326
rect 48412 39976 48464 39982
rect 48412 39918 48464 39924
rect 49056 39976 49108 39982
rect 49056 39918 49108 39924
rect 48424 39642 48452 39918
rect 48596 39840 48648 39846
rect 48596 39782 48648 39788
rect 48964 39840 49016 39846
rect 48964 39782 49016 39788
rect 48608 39642 48636 39782
rect 48412 39636 48464 39642
rect 48412 39578 48464 39584
rect 48596 39636 48648 39642
rect 48596 39578 48648 39584
rect 48320 39092 48372 39098
rect 48320 39034 48372 39040
rect 48332 38962 48360 39034
rect 48320 38956 48372 38962
rect 48320 38898 48372 38904
rect 48228 38412 48280 38418
rect 48228 38354 48280 38360
rect 47860 37868 47912 37874
rect 47860 37810 47912 37816
rect 47860 37732 47912 37738
rect 48240 37720 48268 38354
rect 48332 37890 48360 38898
rect 48424 38894 48452 39578
rect 48976 39098 49004 39782
rect 49160 39681 49188 40718
rect 49146 39672 49202 39681
rect 49146 39607 49202 39616
rect 48964 39092 49016 39098
rect 48964 39034 49016 39040
rect 49344 38962 49372 41074
rect 49516 40996 49568 41002
rect 49516 40938 49568 40944
rect 49608 40996 49660 41002
rect 49608 40938 49660 40944
rect 49424 40928 49476 40934
rect 49424 40870 49476 40876
rect 49436 40662 49464 40870
rect 49424 40656 49476 40662
rect 49424 40598 49476 40604
rect 49528 40118 49556 40938
rect 49620 40186 49648 40938
rect 50160 40928 50212 40934
rect 50632 40905 50660 41074
rect 50160 40870 50212 40876
rect 50618 40896 50674 40905
rect 49976 40656 50028 40662
rect 49976 40598 50028 40604
rect 49608 40180 49660 40186
rect 49608 40122 49660 40128
rect 49516 40112 49568 40118
rect 49516 40054 49568 40060
rect 49988 39982 50016 40598
rect 50172 40526 50200 40870
rect 50618 40831 50674 40840
rect 50632 40644 50660 40831
rect 50712 40656 50764 40662
rect 50632 40616 50712 40644
rect 50712 40598 50764 40604
rect 50160 40520 50212 40526
rect 50160 40462 50212 40468
rect 50712 40520 50764 40526
rect 50712 40462 50764 40468
rect 49976 39976 50028 39982
rect 49976 39918 50028 39924
rect 49792 39908 49844 39914
rect 49792 39850 49844 39856
rect 49608 39568 49660 39574
rect 49660 39516 49740 39522
rect 49608 39510 49740 39516
rect 49620 39494 49740 39510
rect 49516 39432 49568 39438
rect 49516 39374 49568 39380
rect 49332 38956 49384 38962
rect 49332 38898 49384 38904
rect 49528 38894 49556 39374
rect 48412 38888 48464 38894
rect 48412 38830 48464 38836
rect 49516 38888 49568 38894
rect 49516 38830 49568 38836
rect 49712 38826 49740 39494
rect 49804 38962 49832 39850
rect 50160 39840 50212 39846
rect 50160 39782 50212 39788
rect 50172 39438 50200 39782
rect 50526 39672 50582 39681
rect 50526 39607 50528 39616
rect 50580 39607 50582 39616
rect 50528 39578 50580 39584
rect 50620 39500 50672 39506
rect 50620 39442 50672 39448
rect 50160 39432 50212 39438
rect 50160 39374 50212 39380
rect 50528 39432 50580 39438
rect 50528 39374 50580 39380
rect 49792 38956 49844 38962
rect 49792 38898 49844 38904
rect 49700 38820 49752 38826
rect 49700 38762 49752 38768
rect 48964 38752 49016 38758
rect 48964 38694 49016 38700
rect 48976 38486 49004 38694
rect 49712 38486 49740 38762
rect 48964 38480 49016 38486
rect 48964 38422 49016 38428
rect 49700 38480 49752 38486
rect 49700 38422 49752 38428
rect 49976 38276 50028 38282
rect 49976 38218 50028 38224
rect 49988 38010 50016 38218
rect 49976 38004 50028 38010
rect 49976 37946 50028 37952
rect 50066 37904 50122 37913
rect 48332 37862 48452 37890
rect 48320 37732 48372 37738
rect 48240 37692 48320 37720
rect 47860 37674 47912 37680
rect 48320 37674 48372 37680
rect 47584 37664 47636 37670
rect 47584 37606 47636 37612
rect 47492 37460 47544 37466
rect 47492 37402 47544 37408
rect 47596 37398 47624 37606
rect 47872 37466 47900 37674
rect 48424 37670 48452 37862
rect 49700 37868 49752 37874
rect 50172 37874 50200 39374
rect 50344 39024 50396 39030
rect 50344 38966 50396 38972
rect 50356 38554 50384 38966
rect 50540 38894 50568 39374
rect 50632 39030 50660 39442
rect 50620 39024 50672 39030
rect 50620 38966 50672 38972
rect 50528 38888 50580 38894
rect 50528 38830 50580 38836
rect 50344 38548 50396 38554
rect 50344 38490 50396 38496
rect 50066 37839 50122 37848
rect 50160 37868 50212 37874
rect 49700 37810 49752 37816
rect 48412 37664 48464 37670
rect 48412 37606 48464 37612
rect 47860 37460 47912 37466
rect 47860 37402 47912 37408
rect 47584 37392 47636 37398
rect 47584 37334 47636 37340
rect 49712 37262 49740 37810
rect 50080 37466 50108 37839
rect 50160 37810 50212 37816
rect 50068 37460 50120 37466
rect 50068 37402 50120 37408
rect 50080 37330 50108 37402
rect 50068 37324 50120 37330
rect 50068 37266 50120 37272
rect 50540 37262 50568 38830
rect 50724 38826 50752 40462
rect 50908 39846 50936 41482
rect 50998 41372 51306 41381
rect 50998 41370 51004 41372
rect 51060 41370 51084 41372
rect 51140 41370 51164 41372
rect 51220 41370 51244 41372
rect 51300 41370 51306 41372
rect 51060 41318 51062 41370
rect 51242 41318 51244 41370
rect 50998 41316 51004 41318
rect 51060 41316 51084 41318
rect 51140 41316 51164 41318
rect 51220 41316 51244 41318
rect 51300 41316 51306 41318
rect 50998 41307 51306 41316
rect 51080 41064 51132 41070
rect 51080 41006 51132 41012
rect 51172 41064 51224 41070
rect 51172 41006 51224 41012
rect 51092 40594 51120 41006
rect 51184 40730 51212 41006
rect 51368 40934 51396 41618
rect 51356 40928 51408 40934
rect 51356 40870 51408 40876
rect 51172 40724 51224 40730
rect 51172 40666 51224 40672
rect 51080 40588 51132 40594
rect 51080 40530 51132 40536
rect 51368 40458 51396 40870
rect 51460 40730 51488 41686
rect 52288 41274 52316 41958
rect 52472 41750 52500 41958
rect 52460 41744 52512 41750
rect 52460 41686 52512 41692
rect 53208 41274 53236 41958
rect 53472 41812 53524 41818
rect 53472 41754 53524 41760
rect 52276 41268 52328 41274
rect 52276 41210 52328 41216
rect 53196 41268 53248 41274
rect 53196 41210 53248 41216
rect 51918 40828 52226 40837
rect 51918 40826 51924 40828
rect 51980 40826 52004 40828
rect 52060 40826 52084 40828
rect 52140 40826 52164 40828
rect 52220 40826 52226 40828
rect 51980 40774 51982 40826
rect 52162 40774 52164 40826
rect 51918 40772 51924 40774
rect 51980 40772 52004 40774
rect 52060 40772 52084 40774
rect 52140 40772 52164 40774
rect 52220 40772 52226 40774
rect 51918 40763 52226 40772
rect 51448 40724 51500 40730
rect 51448 40666 51500 40672
rect 52288 40594 52316 41210
rect 52552 41200 52604 41206
rect 52552 41142 52604 41148
rect 52368 40928 52420 40934
rect 52368 40870 52420 40876
rect 52380 40730 52408 40870
rect 52368 40724 52420 40730
rect 52368 40666 52420 40672
rect 52276 40588 52328 40594
rect 52276 40530 52328 40536
rect 51816 40520 51868 40526
rect 51816 40462 51868 40468
rect 51356 40452 51408 40458
rect 51356 40394 51408 40400
rect 50998 40284 51306 40293
rect 50998 40282 51004 40284
rect 51060 40282 51084 40284
rect 51140 40282 51164 40284
rect 51220 40282 51244 40284
rect 51300 40282 51306 40284
rect 51060 40230 51062 40282
rect 51242 40230 51244 40282
rect 50998 40228 51004 40230
rect 51060 40228 51084 40230
rect 51140 40228 51164 40230
rect 51220 40228 51244 40230
rect 51300 40228 51306 40230
rect 50998 40219 51306 40228
rect 51828 40186 51856 40462
rect 51816 40180 51868 40186
rect 51816 40122 51868 40128
rect 52460 40044 52512 40050
rect 52460 39986 52512 39992
rect 50896 39840 50948 39846
rect 50896 39782 50948 39788
rect 51918 39740 52226 39749
rect 51918 39738 51924 39740
rect 51980 39738 52004 39740
rect 52060 39738 52084 39740
rect 52140 39738 52164 39740
rect 52220 39738 52226 39740
rect 51980 39686 51982 39738
rect 52162 39686 52164 39738
rect 51918 39684 51924 39686
rect 51980 39684 52004 39686
rect 52060 39684 52084 39686
rect 52140 39684 52164 39686
rect 52220 39684 52226 39686
rect 51918 39675 52226 39684
rect 50804 39500 50856 39506
rect 50804 39442 50856 39448
rect 50816 38962 50844 39442
rect 50998 39196 51306 39205
rect 50998 39194 51004 39196
rect 51060 39194 51084 39196
rect 51140 39194 51164 39196
rect 51220 39194 51244 39196
rect 51300 39194 51306 39196
rect 51060 39142 51062 39194
rect 51242 39142 51244 39194
rect 50998 39140 51004 39142
rect 51060 39140 51084 39142
rect 51140 39140 51164 39142
rect 51220 39140 51244 39142
rect 51300 39140 51306 39142
rect 50998 39131 51306 39140
rect 52472 38962 52500 39986
rect 52564 39506 52592 41142
rect 52828 40928 52880 40934
rect 52828 40870 52880 40876
rect 52840 40526 52868 40870
rect 53484 40594 53512 41754
rect 54036 41206 54064 41958
rect 54128 41546 54156 42638
rect 54208 42220 54260 42226
rect 54208 42162 54260 42168
rect 54116 41540 54168 41546
rect 54116 41482 54168 41488
rect 54024 41200 54076 41206
rect 54024 41142 54076 41148
rect 54220 41138 54248 42162
rect 54484 42084 54536 42090
rect 54484 42026 54536 42032
rect 54496 41206 54524 42026
rect 54852 42016 54904 42022
rect 54852 41958 54904 41964
rect 54864 41206 54892 41958
rect 58348 41812 58400 41818
rect 58348 41754 58400 41760
rect 55128 41676 55180 41682
rect 55128 41618 55180 41624
rect 57704 41676 57756 41682
rect 57704 41618 57756 41624
rect 54944 41540 54996 41546
rect 54944 41482 54996 41488
rect 54484 41200 54536 41206
rect 54484 41142 54536 41148
rect 54852 41200 54904 41206
rect 54852 41142 54904 41148
rect 53656 41132 53708 41138
rect 53656 41074 53708 41080
rect 54208 41132 54260 41138
rect 54208 41074 54260 41080
rect 53472 40588 53524 40594
rect 53472 40530 53524 40536
rect 52828 40520 52880 40526
rect 52828 40462 52880 40468
rect 52840 39914 52868 40462
rect 53564 40384 53616 40390
rect 53668 40338 53696 41074
rect 54220 40526 54248 41074
rect 54208 40520 54260 40526
rect 54208 40462 54260 40468
rect 54496 40390 54524 41142
rect 54864 41018 54892 41142
rect 54772 41002 54892 41018
rect 54760 40996 54892 41002
rect 54812 40990 54892 40996
rect 54760 40938 54812 40944
rect 54576 40520 54628 40526
rect 54576 40462 54628 40468
rect 53616 40332 53696 40338
rect 53564 40326 53696 40332
rect 54484 40384 54536 40390
rect 54484 40326 54536 40332
rect 53576 40310 53696 40326
rect 53668 40050 53696 40310
rect 53656 40044 53708 40050
rect 53656 39986 53708 39992
rect 52828 39908 52880 39914
rect 52828 39850 52880 39856
rect 52552 39500 52604 39506
rect 52552 39442 52604 39448
rect 52736 39296 52788 39302
rect 52736 39238 52788 39244
rect 50804 38956 50856 38962
rect 50804 38898 50856 38904
rect 52460 38956 52512 38962
rect 52460 38898 52512 38904
rect 50712 38820 50764 38826
rect 50712 38762 50764 38768
rect 50816 38418 50844 38898
rect 52276 38888 52328 38894
rect 52276 38830 52328 38836
rect 50988 38752 51040 38758
rect 50988 38694 51040 38700
rect 51000 38554 51028 38694
rect 51918 38652 52226 38661
rect 51918 38650 51924 38652
rect 51980 38650 52004 38652
rect 52060 38650 52084 38652
rect 52140 38650 52164 38652
rect 52220 38650 52226 38652
rect 51980 38598 51982 38650
rect 52162 38598 52164 38650
rect 51918 38596 51924 38598
rect 51980 38596 52004 38598
rect 52060 38596 52084 38598
rect 52140 38596 52164 38598
rect 52220 38596 52226 38598
rect 51918 38587 52226 38596
rect 50988 38548 51040 38554
rect 50988 38490 51040 38496
rect 50804 38412 50856 38418
rect 50804 38354 50856 38360
rect 50896 38344 50948 38350
rect 50896 38286 50948 38292
rect 51724 38344 51776 38350
rect 51724 38286 51776 38292
rect 50620 38208 50672 38214
rect 50620 38150 50672 38156
rect 50632 38010 50660 38150
rect 50620 38004 50672 38010
rect 50620 37946 50672 37952
rect 50712 38004 50764 38010
rect 50712 37946 50764 37952
rect 50724 37466 50752 37946
rect 50908 37466 50936 38286
rect 51632 38208 51684 38214
rect 51632 38150 51684 38156
rect 50998 38108 51306 38117
rect 50998 38106 51004 38108
rect 51060 38106 51084 38108
rect 51140 38106 51164 38108
rect 51220 38106 51244 38108
rect 51300 38106 51306 38108
rect 51060 38054 51062 38106
rect 51242 38054 51244 38106
rect 50998 38052 51004 38054
rect 51060 38052 51084 38054
rect 51140 38052 51164 38054
rect 51220 38052 51244 38054
rect 51300 38052 51306 38054
rect 50998 38043 51306 38052
rect 50712 37460 50764 37466
rect 50712 37402 50764 37408
rect 50896 37460 50948 37466
rect 50896 37402 50948 37408
rect 51644 37398 51672 38150
rect 51736 38010 51764 38286
rect 51724 38004 51776 38010
rect 51724 37946 51776 37952
rect 51724 37664 51776 37670
rect 51724 37606 51776 37612
rect 51816 37664 51868 37670
rect 51816 37606 51868 37612
rect 51736 37398 51764 37606
rect 51632 37392 51684 37398
rect 51632 37334 51684 37340
rect 51724 37392 51776 37398
rect 51724 37334 51776 37340
rect 51828 37330 51856 37606
rect 51918 37564 52226 37573
rect 51918 37562 51924 37564
rect 51980 37562 52004 37564
rect 52060 37562 52084 37564
rect 52140 37562 52164 37564
rect 52220 37562 52226 37564
rect 51980 37510 51982 37562
rect 52162 37510 52164 37562
rect 51918 37508 51924 37510
rect 51980 37508 52004 37510
rect 52060 37508 52084 37510
rect 52140 37508 52164 37510
rect 52220 37508 52226 37510
rect 51918 37499 52226 37508
rect 52288 37398 52316 38830
rect 52748 38826 52776 39238
rect 52840 39001 52868 39850
rect 53668 39658 53696 39986
rect 53748 39976 53800 39982
rect 53748 39918 53800 39924
rect 53576 39630 53696 39658
rect 52826 38992 52882 39001
rect 52826 38927 52882 38936
rect 53472 38956 53524 38962
rect 53472 38898 53524 38904
rect 52736 38820 52788 38826
rect 52736 38762 52788 38768
rect 53484 37806 53512 38898
rect 53472 37800 53524 37806
rect 53472 37742 53524 37748
rect 53196 37732 53248 37738
rect 53196 37674 53248 37680
rect 52276 37392 52328 37398
rect 52276 37334 52328 37340
rect 53208 37330 53236 37674
rect 51816 37324 51868 37330
rect 51816 37266 51868 37272
rect 53196 37324 53248 37330
rect 53196 37266 53248 37272
rect 53576 37262 53604 39630
rect 53760 39574 53788 39918
rect 53748 39568 53800 39574
rect 53748 39510 53800 39516
rect 54496 39522 54524 40326
rect 54588 39642 54616 40462
rect 54956 39642 54984 41482
rect 55036 41132 55088 41138
rect 55036 41074 55088 41080
rect 55048 40934 55076 41074
rect 55036 40928 55088 40934
rect 55036 40870 55088 40876
rect 54576 39636 54628 39642
rect 54576 39578 54628 39584
rect 54944 39636 54996 39642
rect 54944 39578 54996 39584
rect 53656 39500 53708 39506
rect 54496 39494 54616 39522
rect 53656 39442 53708 39448
rect 53668 37330 53696 39442
rect 54588 39438 54616 39494
rect 55048 39438 55076 40870
rect 55140 40730 55168 41618
rect 56140 41608 56192 41614
rect 56140 41550 56192 41556
rect 56508 41608 56560 41614
rect 56508 41550 56560 41556
rect 55680 41472 55732 41478
rect 55680 41414 55732 41420
rect 55692 40934 55720 41414
rect 56152 40934 56180 41550
rect 56416 41472 56468 41478
rect 56416 41414 56468 41420
rect 56428 41070 56456 41414
rect 56416 41064 56468 41070
rect 56416 41006 56468 41012
rect 55220 40928 55272 40934
rect 55220 40870 55272 40876
rect 55680 40928 55732 40934
rect 55680 40870 55732 40876
rect 55772 40928 55824 40934
rect 55772 40870 55824 40876
rect 56140 40928 56192 40934
rect 56140 40870 56192 40876
rect 55128 40724 55180 40730
rect 55128 40666 55180 40672
rect 54484 39432 54536 39438
rect 54484 39374 54536 39380
rect 54576 39432 54628 39438
rect 54576 39374 54628 39380
rect 54852 39432 54904 39438
rect 54852 39374 54904 39380
rect 55036 39432 55088 39438
rect 55036 39374 55088 39380
rect 54208 39364 54260 39370
rect 54208 39306 54260 39312
rect 54220 39098 54248 39306
rect 54496 39098 54524 39374
rect 54208 39092 54260 39098
rect 54208 39034 54260 39040
rect 54484 39092 54536 39098
rect 54484 39034 54536 39040
rect 53840 38888 53892 38894
rect 53840 38830 53892 38836
rect 53852 38486 53880 38830
rect 54116 38752 54168 38758
rect 54116 38694 54168 38700
rect 53840 38480 53892 38486
rect 53840 38422 53892 38428
rect 53852 37942 53880 38422
rect 54128 38350 54156 38694
rect 54116 38344 54168 38350
rect 53944 38304 54116 38332
rect 53840 37936 53892 37942
rect 53840 37878 53892 37884
rect 53944 37738 53972 38304
rect 54116 38286 54168 38292
rect 54220 37738 54248 39034
rect 54588 39030 54616 39374
rect 54576 39024 54628 39030
rect 54576 38966 54628 38972
rect 54392 38344 54444 38350
rect 54392 38286 54444 38292
rect 54404 38010 54432 38286
rect 54392 38004 54444 38010
rect 54392 37946 54444 37952
rect 53932 37732 53984 37738
rect 53932 37674 53984 37680
rect 54208 37732 54260 37738
rect 54208 37674 54260 37680
rect 53656 37324 53708 37330
rect 53656 37266 53708 37272
rect 40868 37256 40920 37262
rect 39684 37194 40080 37210
rect 40868 37198 40920 37204
rect 41236 37256 41288 37262
rect 41236 37198 41288 37204
rect 47124 37256 47176 37262
rect 47124 37198 47176 37204
rect 47308 37256 47360 37262
rect 47308 37198 47360 37204
rect 49700 37256 49752 37262
rect 49700 37198 49752 37204
rect 50528 37256 50580 37262
rect 50528 37198 50580 37204
rect 51448 37256 51500 37262
rect 51448 37198 51500 37204
rect 53564 37256 53616 37262
rect 53564 37198 53616 37204
rect 39672 37188 40092 37194
rect 39724 37182 40040 37188
rect 39672 37130 39724 37136
rect 40040 37130 40092 37136
rect 50998 37020 51306 37029
rect 50998 37018 51004 37020
rect 51060 37018 51084 37020
rect 51140 37018 51164 37020
rect 51220 37018 51244 37020
rect 51300 37018 51306 37020
rect 51060 36966 51062 37018
rect 51242 36966 51244 37018
rect 50998 36964 51004 36966
rect 51060 36964 51084 36966
rect 51140 36964 51164 36966
rect 51220 36964 51244 36966
rect 51300 36964 51306 36966
rect 50998 36955 51306 36964
rect 51460 36922 51488 37198
rect 54588 36922 54616 38966
rect 54864 37874 54892 39374
rect 55140 38894 55168 40666
rect 55232 40662 55260 40870
rect 55220 40656 55272 40662
rect 55220 40598 55272 40604
rect 55784 40526 55812 40870
rect 55772 40520 55824 40526
rect 55772 40462 55824 40468
rect 55680 40044 55732 40050
rect 55680 39986 55732 39992
rect 55312 39908 55364 39914
rect 55312 39850 55364 39856
rect 55220 39840 55272 39846
rect 55220 39782 55272 39788
rect 55232 39302 55260 39782
rect 55324 39642 55352 39850
rect 55312 39636 55364 39642
rect 55312 39578 55364 39584
rect 55220 39296 55272 39302
rect 55220 39238 55272 39244
rect 55232 38962 55260 39238
rect 55692 38962 55720 39986
rect 55784 39846 55812 40462
rect 55772 39840 55824 39846
rect 55772 39782 55824 39788
rect 55956 39636 56008 39642
rect 55956 39578 56008 39584
rect 55220 38956 55272 38962
rect 55220 38898 55272 38904
rect 55680 38956 55732 38962
rect 55680 38898 55732 38904
rect 55968 38894 55996 39578
rect 56520 39574 56548 41550
rect 57716 41274 57744 41618
rect 57796 41472 57848 41478
rect 57796 41414 57848 41420
rect 57704 41268 57756 41274
rect 57704 41210 57756 41216
rect 56692 41132 56744 41138
rect 56692 41074 56744 41080
rect 57060 41132 57112 41138
rect 57060 41074 57112 41080
rect 56600 40996 56652 41002
rect 56600 40938 56652 40944
rect 56612 40186 56640 40938
rect 56704 40730 56732 41074
rect 57072 41002 57100 41074
rect 57612 41064 57664 41070
rect 57612 41006 57664 41012
rect 57060 40996 57112 41002
rect 57060 40938 57112 40944
rect 57520 40996 57572 41002
rect 57520 40938 57572 40944
rect 56692 40724 56744 40730
rect 56692 40666 56744 40672
rect 56704 40390 56732 40666
rect 57072 40633 57100 40938
rect 57152 40928 57204 40934
rect 57152 40870 57204 40876
rect 57058 40624 57114 40633
rect 57058 40559 57114 40568
rect 56692 40384 56744 40390
rect 56692 40326 56744 40332
rect 56600 40180 56652 40186
rect 56600 40122 56652 40128
rect 57164 40118 57192 40870
rect 57532 40730 57560 40938
rect 57520 40724 57572 40730
rect 57520 40666 57572 40672
rect 57532 40186 57560 40666
rect 57624 40610 57652 41006
rect 57716 40730 57744 41210
rect 57704 40724 57756 40730
rect 57704 40666 57756 40672
rect 57808 40610 57836 41414
rect 57624 40582 57836 40610
rect 57520 40180 57572 40186
rect 57520 40122 57572 40128
rect 57152 40112 57204 40118
rect 57152 40054 57204 40060
rect 57336 39908 57388 39914
rect 57336 39850 57388 39856
rect 57244 39840 57296 39846
rect 57244 39782 57296 39788
rect 57256 39574 57284 39782
rect 56508 39568 56560 39574
rect 56508 39510 56560 39516
rect 57244 39568 57296 39574
rect 57244 39510 57296 39516
rect 56140 39296 56192 39302
rect 56140 39238 56192 39244
rect 56152 38894 56180 39238
rect 56520 38962 56548 39510
rect 57348 39438 57376 39850
rect 57152 39432 57204 39438
rect 57152 39374 57204 39380
rect 57336 39432 57388 39438
rect 57336 39374 57388 39380
rect 56508 38956 56560 38962
rect 56508 38898 56560 38904
rect 55128 38888 55180 38894
rect 55128 38830 55180 38836
rect 55956 38888 56008 38894
rect 55956 38830 56008 38836
rect 56140 38888 56192 38894
rect 56140 38830 56192 38836
rect 55128 38752 55180 38758
rect 55128 38694 55180 38700
rect 55772 38752 55824 38758
rect 55772 38694 55824 38700
rect 54852 37868 54904 37874
rect 54852 37810 54904 37816
rect 54864 37262 54892 37810
rect 55140 37738 55168 38694
rect 55784 38486 55812 38694
rect 55968 38486 55996 38830
rect 56232 38752 56284 38758
rect 56232 38694 56284 38700
rect 55772 38480 55824 38486
rect 55772 38422 55824 38428
rect 55956 38480 56008 38486
rect 55956 38422 56008 38428
rect 55220 38344 55272 38350
rect 55220 38286 55272 38292
rect 55232 37806 55260 38286
rect 55220 37800 55272 37806
rect 55220 37742 55272 37748
rect 55402 37768 55458 37777
rect 55128 37732 55180 37738
rect 55128 37674 55180 37680
rect 55232 37398 55260 37742
rect 55402 37703 55404 37712
rect 55456 37703 55458 37712
rect 55862 37768 55918 37777
rect 55968 37738 55996 38422
rect 56244 38010 56272 38694
rect 56784 38276 56836 38282
rect 56784 38218 56836 38224
rect 56232 38004 56284 38010
rect 56232 37946 56284 37952
rect 56600 37936 56652 37942
rect 56600 37878 56652 37884
rect 55862 37703 55864 37712
rect 55404 37674 55456 37680
rect 55916 37703 55918 37712
rect 55956 37732 56008 37738
rect 55864 37674 55916 37680
rect 55956 37674 56008 37680
rect 55220 37392 55272 37398
rect 55220 37334 55272 37340
rect 56416 37392 56468 37398
rect 56416 37334 56468 37340
rect 54852 37256 54904 37262
rect 54852 37198 54904 37204
rect 56428 37126 56456 37334
rect 56612 37194 56640 37878
rect 56796 37466 56824 38218
rect 57164 38214 57192 39374
rect 57152 38208 57204 38214
rect 57152 38150 57204 38156
rect 57336 37732 57388 37738
rect 57336 37674 57388 37680
rect 57348 37466 57376 37674
rect 56784 37460 56836 37466
rect 56784 37402 56836 37408
rect 57336 37460 57388 37466
rect 57336 37402 57388 37408
rect 57624 37194 57652 40582
rect 57704 39976 57756 39982
rect 57702 39944 57704 39953
rect 57756 39944 57758 39953
rect 57702 39879 57758 39888
rect 57716 39438 57744 39879
rect 58072 39840 58124 39846
rect 58072 39782 58124 39788
rect 57704 39432 57756 39438
rect 57704 39374 57756 39380
rect 57796 39296 57848 39302
rect 57796 39238 57848 39244
rect 57808 38350 57836 39238
rect 58084 39098 58112 39782
rect 58072 39092 58124 39098
rect 58072 39034 58124 39040
rect 57980 38956 58032 38962
rect 57980 38898 58032 38904
rect 57796 38344 57848 38350
rect 57848 38304 57928 38332
rect 57796 38286 57848 38292
rect 57704 38208 57756 38214
rect 57704 38150 57756 38156
rect 57716 37466 57744 38150
rect 57900 38010 57928 38304
rect 57888 38004 57940 38010
rect 57888 37946 57940 37952
rect 57900 37874 57928 37946
rect 57992 37874 58020 38898
rect 58360 38826 58388 41754
rect 58716 40112 58768 40118
rect 58716 40054 58768 40060
rect 58440 39840 58492 39846
rect 58440 39782 58492 39788
rect 58452 39642 58480 39782
rect 58440 39636 58492 39642
rect 58440 39578 58492 39584
rect 58348 38820 58400 38826
rect 58348 38762 58400 38768
rect 58360 38486 58388 38762
rect 58348 38480 58400 38486
rect 58348 38422 58400 38428
rect 58164 38344 58216 38350
rect 58164 38286 58216 38292
rect 58360 38332 58388 38422
rect 58440 38344 58492 38350
rect 58360 38304 58440 38332
rect 57888 37868 57940 37874
rect 57888 37810 57940 37816
rect 57980 37868 58032 37874
rect 57980 37810 58032 37816
rect 57796 37664 57848 37670
rect 57796 37606 57848 37612
rect 57808 37466 57836 37606
rect 58176 37466 58204 38286
rect 58360 37806 58388 38304
rect 58440 38286 58492 38292
rect 58440 37936 58492 37942
rect 58440 37878 58492 37884
rect 58348 37800 58400 37806
rect 58348 37742 58400 37748
rect 58452 37754 58480 37878
rect 58452 37726 58664 37754
rect 58532 37664 58584 37670
rect 58532 37606 58584 37612
rect 58544 37466 58572 37606
rect 58636 37466 58664 37726
rect 57704 37460 57756 37466
rect 57704 37402 57756 37408
rect 57796 37460 57848 37466
rect 57796 37402 57848 37408
rect 58164 37460 58216 37466
rect 58164 37402 58216 37408
rect 58532 37460 58584 37466
rect 58532 37402 58584 37408
rect 58624 37460 58676 37466
rect 58624 37402 58676 37408
rect 57808 37330 57836 37402
rect 57796 37324 57848 37330
rect 57796 37266 57848 37272
rect 58728 37262 58756 40054
rect 58808 39908 58860 39914
rect 58808 39850 58860 39856
rect 58820 39370 58848 39850
rect 58900 39840 58952 39846
rect 58900 39782 58952 39788
rect 58808 39364 58860 39370
rect 58808 39306 58860 39312
rect 58820 39098 58848 39306
rect 58912 39098 58940 39782
rect 59268 39432 59320 39438
rect 59268 39374 59320 39380
rect 58808 39092 58860 39098
rect 58808 39034 58860 39040
rect 58900 39092 58952 39098
rect 58900 39034 58952 39040
rect 59280 38894 59308 39374
rect 59452 38956 59504 38962
rect 59452 38898 59504 38904
rect 59268 38888 59320 38894
rect 59268 38830 59320 38836
rect 59268 38752 59320 38758
rect 59268 38694 59320 38700
rect 59280 38350 59308 38694
rect 59268 38344 59320 38350
rect 59268 38286 59320 38292
rect 59280 37466 59308 38286
rect 59268 37460 59320 37466
rect 59268 37402 59320 37408
rect 58716 37256 58768 37262
rect 58716 37198 58768 37204
rect 59464 37194 59492 38898
rect 60016 37806 60044 42706
rect 60738 42664 60794 42673
rect 60738 42599 60794 42608
rect 60648 40724 60700 40730
rect 60648 40666 60700 40672
rect 60660 39930 60688 40666
rect 60752 40225 60780 42599
rect 65800 42560 65852 42566
rect 65800 42502 65852 42508
rect 63040 42152 63092 42158
rect 63040 42094 63092 42100
rect 62854 41032 62910 41041
rect 62854 40967 62910 40976
rect 60738 40216 60794 40225
rect 60738 40151 60794 40160
rect 60660 39902 60780 39930
rect 60752 38486 60780 39902
rect 60740 38480 60792 38486
rect 60740 38422 60792 38428
rect 62488 38480 62540 38486
rect 62488 38422 62540 38428
rect 60004 37800 60056 37806
rect 60004 37742 60056 37748
rect 59820 37732 59872 37738
rect 59820 37674 59872 37680
rect 59832 37466 59860 37674
rect 60280 37664 60332 37670
rect 60280 37606 60332 37612
rect 60292 37466 60320 37606
rect 59728 37460 59780 37466
rect 59728 37402 59780 37408
rect 59820 37460 59872 37466
rect 59820 37402 59872 37408
rect 60280 37460 60332 37466
rect 60280 37402 60332 37408
rect 59740 37346 59768 37402
rect 62026 37360 62082 37369
rect 59740 37330 59952 37346
rect 59740 37324 59964 37330
rect 59740 37318 59912 37324
rect 62026 37295 62082 37304
rect 59912 37266 59964 37272
rect 60464 37256 60516 37262
rect 60464 37198 60516 37204
rect 56600 37188 56652 37194
rect 56600 37130 56652 37136
rect 57612 37188 57664 37194
rect 57612 37130 57664 37136
rect 59452 37188 59504 37194
rect 59452 37130 59504 37136
rect 56416 37120 56468 37126
rect 56416 37062 56468 37068
rect 51448 36916 51500 36922
rect 51448 36858 51500 36864
rect 54576 36916 54628 36922
rect 54576 36858 54628 36864
rect 38568 36780 38620 36786
rect 38568 36722 38620 36728
rect 38752 36780 38804 36786
rect 38752 36722 38804 36728
rect 34428 36644 34480 36650
rect 34428 36586 34480 36592
rect 37648 36644 37700 36650
rect 37648 36586 37700 36592
rect 34440 36145 34468 36586
rect 37280 36508 37332 36514
rect 37280 36450 37332 36456
rect 37292 36281 37320 36450
rect 37278 36272 37334 36281
rect 37278 36207 37334 36216
rect 34426 36136 34482 36145
rect 34426 36071 34482 36080
rect 36544 35896 36596 35902
rect 34518 35864 34574 35873
rect 34164 35822 34518 35850
rect 33046 35799 33102 35808
rect 38580 35873 38608 36722
rect 38660 36712 38712 36718
rect 38660 36654 38712 36660
rect 36544 35838 36596 35844
rect 38566 35864 38622 35873
rect 34518 35799 34574 35808
rect 36556 35737 36584 35838
rect 38566 35799 38622 35808
rect 38672 35737 38700 36654
rect 42708 36372 42760 36378
rect 42708 36314 42760 36320
rect 42616 36236 42668 36242
rect 42616 36178 42668 36184
rect 30286 35728 30342 35737
rect 30470 35728 30526 35737
rect 30286 35663 30342 35672
rect 30392 35686 30470 35714
rect 30392 35578 30420 35686
rect 30470 35663 30526 35672
rect 36542 35728 36598 35737
rect 36542 35663 36598 35672
rect 38658 35728 38714 35737
rect 42628 35698 42656 36178
rect 42720 35873 42748 36314
rect 42706 35864 42762 35873
rect 42706 35799 42762 35808
rect 56428 35737 56456 37062
rect 60476 36854 60504 37198
rect 60464 36848 60516 36854
rect 60464 36790 60516 36796
rect 60832 36576 60884 36582
rect 60832 36518 60884 36524
rect 59360 36236 59412 36242
rect 59360 36178 59412 36184
rect 59372 35766 59400 36178
rect 59360 35760 59412 35766
rect 56414 35728 56470 35737
rect 38658 35663 38714 35672
rect 42616 35692 42668 35698
rect 59360 35702 59412 35708
rect 56414 35663 56470 35672
rect 42616 35634 42668 35640
rect 29932 35550 30420 35578
rect 60844 35562 60872 36518
rect 62040 35630 62068 37295
rect 62120 36168 62172 36174
rect 62120 36110 62172 36116
rect 62132 36009 62160 36110
rect 62118 36000 62174 36009
rect 62118 35935 62174 35944
rect 62028 35624 62080 35630
rect 62028 35566 62080 35572
rect 60832 35556 60884 35562
rect 60832 35498 60884 35504
rect 62500 34950 62528 38422
rect 62764 37392 62816 37398
rect 62764 37334 62816 37340
rect 62578 36272 62634 36281
rect 62578 36207 62634 36216
rect 62488 34944 62540 34950
rect 62488 34886 62540 34892
rect 62592 31090 62620 36207
rect 62670 36136 62726 36145
rect 62670 36071 62726 36080
rect 62684 31249 62712 36071
rect 62670 31240 62726 31249
rect 62670 31175 62726 31184
rect 62592 31062 62712 31090
rect 62580 31000 62632 31006
rect 62580 30942 62632 30948
rect 49240 2032 49292 2038
rect 49240 1974 49292 1980
rect 48964 1964 49016 1970
rect 48964 1906 49016 1912
rect 48976 1873 49004 1906
rect 49252 1873 49280 1974
rect 49700 1896 49752 1902
rect 48962 1864 49018 1873
rect 48962 1799 49018 1808
rect 49238 1864 49294 1873
rect 49238 1799 49294 1808
rect 49698 1864 49700 1873
rect 49752 1864 49754 1873
rect 49698 1799 49754 1808
rect 62592 1329 62620 30942
rect 62684 1970 62712 31062
rect 62776 23662 62804 37334
rect 62868 33250 62896 40967
rect 62948 37120 63000 37126
rect 62948 37062 63000 37068
rect 62856 33244 62908 33250
rect 62856 33186 62908 33192
rect 62856 27600 62908 27606
rect 62856 27542 62908 27548
rect 62764 23656 62816 23662
rect 62764 23598 62816 23604
rect 62764 15360 62816 15366
rect 62764 15302 62816 15308
rect 62776 2038 62804 15302
rect 62764 2032 62816 2038
rect 62764 1974 62816 1980
rect 62672 1964 62724 1970
rect 62672 1906 62724 1912
rect 62868 1601 62896 27542
rect 62960 14822 62988 37062
rect 63052 23798 63080 42094
rect 64880 40928 64932 40934
rect 64880 40870 64932 40876
rect 63684 38820 63736 38826
rect 63684 38762 63736 38768
rect 63222 38312 63278 38321
rect 63222 38247 63278 38256
rect 63132 37868 63184 37874
rect 63132 37810 63184 37816
rect 63144 37330 63172 37810
rect 63132 37324 63184 37330
rect 63132 37266 63184 37272
rect 63132 36100 63184 36106
rect 63132 36042 63184 36048
rect 63040 23792 63092 23798
rect 63040 23734 63092 23740
rect 63144 23050 63172 36042
rect 63236 31006 63264 38247
rect 63316 38208 63368 38214
rect 63316 38150 63368 38156
rect 63328 34746 63356 38150
rect 63696 37874 63724 38762
rect 63776 38548 63828 38554
rect 63776 38490 63828 38496
rect 63788 37874 63816 38490
rect 63868 38004 63920 38010
rect 63868 37946 63920 37952
rect 63684 37868 63736 37874
rect 63684 37810 63736 37816
rect 63776 37868 63828 37874
rect 63776 37810 63828 37816
rect 63408 37256 63460 37262
rect 63408 37198 63460 37204
rect 63420 36922 63448 37198
rect 63408 36916 63460 36922
rect 63408 36858 63460 36864
rect 63500 36644 63552 36650
rect 63500 36586 63552 36592
rect 63512 35894 63540 36586
rect 63592 36304 63644 36310
rect 63590 36272 63592 36281
rect 63644 36272 63646 36281
rect 63590 36207 63646 36216
rect 63512 35866 63632 35894
rect 63500 35556 63552 35562
rect 63500 35498 63552 35504
rect 63512 34785 63540 35498
rect 63498 34776 63554 34785
rect 63316 34740 63368 34746
rect 63498 34711 63554 34720
rect 63316 34682 63368 34688
rect 63408 33244 63460 33250
rect 63408 33186 63460 33192
rect 63420 31770 63448 33186
rect 63420 31742 63540 31770
rect 63224 31000 63276 31006
rect 63224 30942 63276 30948
rect 63512 27606 63540 31742
rect 63500 27600 63552 27606
rect 63500 27542 63552 27548
rect 63604 27418 63632 35866
rect 63696 35698 63724 37810
rect 63776 36780 63828 36786
rect 63776 36722 63828 36728
rect 63684 35692 63736 35698
rect 63684 35634 63736 35640
rect 63682 34640 63738 34649
rect 63682 34575 63738 34584
rect 63696 31890 63724 34575
rect 63684 31884 63736 31890
rect 63684 31826 63736 31832
rect 63512 27390 63632 27418
rect 63408 23520 63460 23526
rect 63408 23462 63460 23468
rect 63132 23044 63184 23050
rect 63132 22986 63184 22992
rect 63316 21480 63368 21486
rect 63316 21422 63368 21428
rect 63328 16454 63356 21422
rect 63316 16448 63368 16454
rect 63316 16390 63368 16396
rect 62948 14816 63000 14822
rect 62948 14758 63000 14764
rect 63040 13864 63092 13870
rect 63040 13806 63092 13812
rect 63052 1902 63080 13806
rect 63420 4282 63448 23462
rect 63408 4276 63460 4282
rect 63408 4218 63460 4224
rect 63040 1896 63092 1902
rect 63512 1873 63540 27390
rect 63788 27282 63816 36722
rect 63880 36174 63908 37946
rect 64236 37664 64288 37670
rect 64236 37606 64288 37612
rect 64248 36786 64276 37606
rect 64788 37120 64840 37126
rect 64788 37062 64840 37068
rect 64338 37020 64646 37029
rect 64338 37018 64344 37020
rect 64400 37018 64424 37020
rect 64480 37018 64504 37020
rect 64560 37018 64584 37020
rect 64640 37018 64646 37020
rect 64400 36966 64402 37018
rect 64582 36966 64584 37018
rect 64338 36964 64344 36966
rect 64400 36964 64424 36966
rect 64480 36964 64504 36966
rect 64560 36964 64584 36966
rect 64640 36964 64646 36966
rect 64338 36955 64646 36964
rect 64800 36854 64828 37062
rect 64788 36848 64840 36854
rect 64788 36790 64840 36796
rect 64236 36780 64288 36786
rect 64236 36722 64288 36728
rect 64696 36780 64748 36786
rect 64696 36722 64748 36728
rect 63868 36168 63920 36174
rect 63868 36110 63920 36116
rect 64236 36168 64288 36174
rect 64236 36110 64288 36116
rect 63880 34542 63908 36110
rect 64248 35834 64276 36110
rect 64338 35932 64646 35941
rect 64338 35930 64344 35932
rect 64400 35930 64424 35932
rect 64480 35930 64504 35932
rect 64560 35930 64584 35932
rect 64640 35930 64646 35932
rect 64400 35878 64402 35930
rect 64582 35878 64584 35930
rect 64338 35876 64344 35878
rect 64400 35876 64424 35878
rect 64480 35876 64504 35878
rect 64560 35876 64584 35878
rect 64640 35876 64646 35878
rect 64338 35867 64646 35876
rect 64236 35828 64288 35834
rect 64236 35770 64288 35776
rect 63958 35728 64014 35737
rect 63958 35663 64014 35672
rect 63868 34536 63920 34542
rect 63868 34478 63920 34484
rect 63880 32026 63908 34478
rect 63972 32910 64000 35663
rect 64236 35488 64288 35494
rect 64236 35430 64288 35436
rect 64052 34944 64104 34950
rect 64052 34886 64104 34892
rect 64064 34082 64092 34886
rect 64144 34468 64196 34474
rect 64144 34410 64196 34416
rect 64156 34202 64184 34410
rect 64144 34196 64196 34202
rect 64144 34138 64196 34144
rect 64064 34054 64184 34082
rect 63960 32904 64012 32910
rect 63960 32846 64012 32852
rect 63868 32020 63920 32026
rect 63868 31962 63920 31968
rect 63868 31884 63920 31890
rect 63868 31826 63920 31832
rect 63604 27254 63816 27282
rect 63604 13870 63632 27254
rect 63880 27044 63908 31826
rect 63972 30802 64000 32846
rect 64052 32020 64104 32026
rect 64052 31962 64104 31968
rect 63960 30796 64012 30802
rect 63960 30738 64012 30744
rect 64064 29170 64092 31962
rect 64052 29164 64104 29170
rect 64052 29106 64104 29112
rect 64156 29050 64184 34054
rect 63696 27016 63908 27044
rect 63972 29022 64184 29050
rect 63696 23526 63724 27016
rect 63972 26234 64000 29022
rect 64052 26376 64104 26382
rect 64052 26318 64104 26324
rect 63788 26206 64000 26234
rect 63684 23520 63736 23526
rect 63684 23462 63736 23468
rect 63684 14816 63736 14822
rect 63684 14758 63736 14764
rect 63592 13864 63644 13870
rect 63592 13806 63644 13812
rect 63696 11286 63724 14758
rect 63684 11280 63736 11286
rect 63684 11222 63736 11228
rect 63788 6866 63816 26206
rect 63960 25356 64012 25362
rect 63960 25298 64012 25304
rect 63972 24614 64000 25298
rect 63960 24608 64012 24614
rect 63960 24550 64012 24556
rect 63972 24206 64000 24550
rect 63960 24200 64012 24206
rect 63960 24142 64012 24148
rect 63868 23792 63920 23798
rect 63868 23734 63920 23740
rect 63880 21486 63908 23734
rect 63972 22030 64000 24142
rect 64064 23526 64092 26318
rect 64248 26234 64276 35430
rect 64338 34844 64646 34853
rect 64338 34842 64344 34844
rect 64400 34842 64424 34844
rect 64480 34842 64504 34844
rect 64560 34842 64584 34844
rect 64640 34842 64646 34844
rect 64400 34790 64402 34842
rect 64582 34790 64584 34842
rect 64338 34788 64344 34790
rect 64400 34788 64424 34790
rect 64480 34788 64504 34790
rect 64560 34788 64584 34790
rect 64640 34788 64646 34790
rect 64338 34779 64646 34788
rect 64708 33998 64736 36722
rect 64788 36032 64840 36038
rect 64788 35974 64840 35980
rect 64696 33992 64748 33998
rect 64696 33934 64748 33940
rect 64696 33856 64748 33862
rect 64696 33798 64748 33804
rect 64338 33756 64646 33765
rect 64338 33754 64344 33756
rect 64400 33754 64424 33756
rect 64480 33754 64504 33756
rect 64560 33754 64584 33756
rect 64640 33754 64646 33756
rect 64400 33702 64402 33754
rect 64582 33702 64584 33754
rect 64338 33700 64344 33702
rect 64400 33700 64424 33702
rect 64480 33700 64504 33702
rect 64560 33700 64584 33702
rect 64640 33700 64646 33702
rect 64338 33691 64646 33700
rect 64338 32668 64646 32677
rect 64338 32666 64344 32668
rect 64400 32666 64424 32668
rect 64480 32666 64504 32668
rect 64560 32666 64584 32668
rect 64640 32666 64646 32668
rect 64400 32614 64402 32666
rect 64582 32614 64584 32666
rect 64338 32612 64344 32614
rect 64400 32612 64424 32614
rect 64480 32612 64504 32614
rect 64560 32612 64584 32614
rect 64640 32612 64646 32614
rect 64338 32603 64646 32612
rect 64708 32570 64736 33798
rect 64800 33522 64828 35974
rect 64892 35894 64920 40870
rect 64972 38412 65024 38418
rect 64972 38354 65024 38360
rect 64984 37398 65012 38354
rect 65258 37564 65566 37573
rect 65258 37562 65264 37564
rect 65320 37562 65344 37564
rect 65400 37562 65424 37564
rect 65480 37562 65504 37564
rect 65560 37562 65566 37564
rect 65320 37510 65322 37562
rect 65502 37510 65504 37562
rect 65258 37508 65264 37510
rect 65320 37508 65344 37510
rect 65400 37508 65424 37510
rect 65480 37508 65504 37510
rect 65560 37508 65566 37510
rect 65258 37499 65566 37508
rect 65156 37460 65208 37466
rect 65156 37402 65208 37408
rect 64972 37392 65024 37398
rect 64972 37334 65024 37340
rect 65168 37330 65196 37402
rect 65708 37392 65760 37398
rect 65708 37334 65760 37340
rect 65156 37324 65208 37330
rect 65156 37266 65208 37272
rect 64972 37120 65024 37126
rect 64972 37062 65024 37068
rect 64984 36650 65012 37062
rect 64972 36644 65024 36650
rect 64972 36586 65024 36592
rect 65064 36576 65116 36582
rect 65064 36518 65116 36524
rect 64892 35866 65012 35894
rect 64788 33516 64840 33522
rect 64788 33458 64840 33464
rect 64880 32904 64932 32910
rect 64880 32846 64932 32852
rect 64892 32570 64920 32846
rect 64696 32564 64748 32570
rect 64696 32506 64748 32512
rect 64880 32564 64932 32570
rect 64880 32506 64932 32512
rect 64880 32292 64932 32298
rect 64880 32234 64932 32240
rect 64892 31890 64920 32234
rect 64984 31958 65012 35866
rect 65076 35630 65104 36518
rect 65168 35698 65196 37266
rect 65258 36476 65566 36485
rect 65258 36474 65264 36476
rect 65320 36474 65344 36476
rect 65400 36474 65424 36476
rect 65480 36474 65504 36476
rect 65560 36474 65566 36476
rect 65320 36422 65322 36474
rect 65502 36422 65504 36474
rect 65258 36420 65264 36422
rect 65320 36420 65344 36422
rect 65400 36420 65424 36422
rect 65480 36420 65504 36422
rect 65560 36420 65566 36422
rect 65258 36411 65566 36420
rect 65616 36372 65668 36378
rect 65616 36314 65668 36320
rect 65432 36304 65484 36310
rect 65432 36246 65484 36252
rect 65156 35692 65208 35698
rect 65156 35634 65208 35640
rect 65064 35624 65116 35630
rect 65444 35578 65472 36246
rect 65064 35566 65116 35572
rect 65168 35550 65472 35578
rect 65168 34474 65196 35550
rect 65258 35388 65566 35397
rect 65258 35386 65264 35388
rect 65320 35386 65344 35388
rect 65400 35386 65424 35388
rect 65480 35386 65504 35388
rect 65560 35386 65566 35388
rect 65320 35334 65322 35386
rect 65502 35334 65504 35386
rect 65258 35332 65264 35334
rect 65320 35332 65344 35334
rect 65400 35332 65424 35334
rect 65480 35332 65504 35334
rect 65560 35332 65566 35334
rect 65258 35323 65566 35332
rect 65628 34950 65656 36314
rect 65720 36310 65748 37334
rect 65708 36304 65760 36310
rect 65708 36246 65760 36252
rect 65708 35760 65760 35766
rect 65708 35702 65760 35708
rect 65616 34944 65668 34950
rect 65616 34886 65668 34892
rect 65616 34740 65668 34746
rect 65616 34682 65668 34688
rect 65156 34468 65208 34474
rect 65156 34410 65208 34416
rect 65258 34300 65566 34309
rect 65258 34298 65264 34300
rect 65320 34298 65344 34300
rect 65400 34298 65424 34300
rect 65480 34298 65504 34300
rect 65560 34298 65566 34300
rect 65320 34246 65322 34298
rect 65502 34246 65504 34298
rect 65258 34244 65264 34246
rect 65320 34244 65344 34246
rect 65400 34244 65424 34246
rect 65480 34244 65504 34246
rect 65560 34244 65566 34246
rect 65258 34235 65566 34244
rect 65628 34066 65656 34682
rect 65616 34060 65668 34066
rect 65616 34002 65668 34008
rect 65064 33516 65116 33522
rect 65064 33458 65116 33464
rect 64972 31952 65024 31958
rect 64972 31894 65024 31900
rect 64880 31884 64932 31890
rect 64880 31826 64932 31832
rect 64338 31580 64646 31589
rect 64338 31578 64344 31580
rect 64400 31578 64424 31580
rect 64480 31578 64504 31580
rect 64560 31578 64584 31580
rect 64640 31578 64646 31580
rect 64400 31526 64402 31578
rect 64582 31526 64584 31578
rect 64338 31524 64344 31526
rect 64400 31524 64424 31526
rect 64480 31524 64504 31526
rect 64560 31524 64584 31526
rect 64640 31524 64646 31526
rect 64338 31515 64646 31524
rect 64880 31340 64932 31346
rect 64880 31282 64932 31288
rect 64696 30728 64748 30734
rect 64696 30670 64748 30676
rect 64338 30492 64646 30501
rect 64338 30490 64344 30492
rect 64400 30490 64424 30492
rect 64480 30490 64504 30492
rect 64560 30490 64584 30492
rect 64640 30490 64646 30492
rect 64400 30438 64402 30490
rect 64582 30438 64584 30490
rect 64338 30436 64344 30438
rect 64400 30436 64424 30438
rect 64480 30436 64504 30438
rect 64560 30436 64584 30438
rect 64640 30436 64646 30438
rect 64338 30427 64646 30436
rect 64708 30394 64736 30670
rect 64696 30388 64748 30394
rect 64696 30330 64748 30336
rect 64696 29504 64748 29510
rect 64696 29446 64748 29452
rect 64338 29404 64646 29413
rect 64338 29402 64344 29404
rect 64400 29402 64424 29404
rect 64480 29402 64504 29404
rect 64560 29402 64584 29404
rect 64640 29402 64646 29404
rect 64400 29350 64402 29402
rect 64582 29350 64584 29402
rect 64338 29348 64344 29350
rect 64400 29348 64424 29350
rect 64480 29348 64504 29350
rect 64560 29348 64584 29350
rect 64640 29348 64646 29350
rect 64338 29339 64646 29348
rect 64708 29170 64736 29446
rect 64696 29164 64748 29170
rect 64696 29106 64748 29112
rect 64892 28914 64920 31282
rect 64984 29073 65012 31894
rect 65076 31498 65104 33458
rect 65628 33454 65656 34002
rect 65616 33448 65668 33454
rect 65616 33390 65668 33396
rect 65156 33312 65208 33318
rect 65156 33254 65208 33260
rect 65616 33312 65668 33318
rect 65616 33254 65668 33260
rect 65168 32434 65196 33254
rect 65258 33212 65566 33221
rect 65258 33210 65264 33212
rect 65320 33210 65344 33212
rect 65400 33210 65424 33212
rect 65480 33210 65504 33212
rect 65560 33210 65566 33212
rect 65320 33158 65322 33210
rect 65502 33158 65504 33210
rect 65258 33156 65264 33158
rect 65320 33156 65344 33158
rect 65400 33156 65424 33158
rect 65480 33156 65504 33158
rect 65560 33156 65566 33158
rect 65258 33147 65566 33156
rect 65248 32768 65300 32774
rect 65248 32710 65300 32716
rect 65156 32428 65208 32434
rect 65156 32370 65208 32376
rect 65260 32366 65288 32710
rect 65628 32366 65656 33254
rect 65248 32360 65300 32366
rect 65248 32302 65300 32308
rect 65616 32360 65668 32366
rect 65616 32302 65668 32308
rect 65720 32298 65748 35702
rect 65812 35086 65840 42502
rect 66076 41064 66128 41070
rect 66076 41006 66128 41012
rect 65984 37732 66036 37738
rect 65984 37674 66036 37680
rect 65892 36848 65944 36854
rect 65892 36790 65944 36796
rect 65904 35850 65932 36790
rect 65996 36786 66024 37674
rect 65984 36780 66036 36786
rect 65984 36722 66036 36728
rect 65996 36378 66024 36722
rect 65984 36372 66036 36378
rect 65984 36314 66036 36320
rect 65904 35822 66024 35850
rect 65892 35692 65944 35698
rect 65892 35634 65944 35640
rect 65800 35080 65852 35086
rect 65800 35022 65852 35028
rect 65800 34944 65852 34950
rect 65800 34886 65852 34892
rect 65708 32292 65760 32298
rect 65708 32234 65760 32240
rect 65616 32224 65668 32230
rect 65616 32166 65668 32172
rect 65258 32124 65566 32133
rect 65258 32122 65264 32124
rect 65320 32122 65344 32124
rect 65400 32122 65424 32124
rect 65480 32122 65504 32124
rect 65560 32122 65566 32124
rect 65320 32070 65322 32122
rect 65502 32070 65504 32122
rect 65258 32068 65264 32070
rect 65320 32068 65344 32070
rect 65400 32068 65424 32070
rect 65480 32068 65504 32070
rect 65560 32068 65566 32070
rect 65258 32059 65566 32068
rect 65076 31470 65196 31498
rect 65064 31408 65116 31414
rect 65064 31350 65116 31356
rect 65076 30258 65104 31350
rect 65064 30252 65116 30258
rect 65064 30194 65116 30200
rect 65064 29776 65116 29782
rect 65064 29718 65116 29724
rect 64970 29064 65026 29073
rect 64970 28999 65026 29008
rect 64892 28886 65012 28914
rect 64878 28792 64934 28801
rect 64878 28727 64934 28736
rect 64338 28316 64646 28325
rect 64338 28314 64344 28316
rect 64400 28314 64424 28316
rect 64480 28314 64504 28316
rect 64560 28314 64584 28316
rect 64640 28314 64646 28316
rect 64400 28262 64402 28314
rect 64582 28262 64584 28314
rect 64338 28260 64344 28262
rect 64400 28260 64424 28262
rect 64480 28260 64504 28262
rect 64560 28260 64584 28262
rect 64640 28260 64646 28262
rect 64338 28251 64646 28260
rect 64338 27228 64646 27237
rect 64338 27226 64344 27228
rect 64400 27226 64424 27228
rect 64480 27226 64504 27228
rect 64560 27226 64584 27228
rect 64640 27226 64646 27228
rect 64400 27174 64402 27226
rect 64582 27174 64584 27226
rect 64338 27172 64344 27174
rect 64400 27172 64424 27174
rect 64480 27172 64504 27174
rect 64560 27172 64584 27174
rect 64640 27172 64646 27174
rect 64338 27163 64646 27172
rect 64696 26376 64748 26382
rect 64696 26318 64748 26324
rect 64156 26206 64276 26234
rect 64052 23520 64104 23526
rect 64052 23462 64104 23468
rect 64064 23186 64092 23462
rect 64052 23180 64104 23186
rect 64052 23122 64104 23128
rect 63960 22024 64012 22030
rect 63960 21966 64012 21972
rect 63868 21480 63920 21486
rect 63868 21422 63920 21428
rect 63972 16574 64000 21966
rect 64064 19922 64092 23122
rect 64156 20754 64184 26206
rect 64338 26140 64646 26149
rect 64338 26138 64344 26140
rect 64400 26138 64424 26140
rect 64480 26138 64504 26140
rect 64560 26138 64584 26140
rect 64640 26138 64646 26140
rect 64400 26086 64402 26138
rect 64582 26086 64584 26138
rect 64338 26084 64344 26086
rect 64400 26084 64424 26086
rect 64480 26084 64504 26086
rect 64560 26084 64584 26086
rect 64640 26084 64646 26086
rect 64338 26075 64646 26084
rect 64708 26042 64736 26318
rect 64696 26036 64748 26042
rect 64696 25978 64748 25984
rect 64236 25152 64288 25158
rect 64236 25094 64288 25100
rect 64248 24342 64276 25094
rect 64338 25052 64646 25061
rect 64338 25050 64344 25052
rect 64400 25050 64424 25052
rect 64480 25050 64504 25052
rect 64560 25050 64584 25052
rect 64640 25050 64646 25052
rect 64400 24998 64402 25050
rect 64582 24998 64584 25050
rect 64338 24996 64344 24998
rect 64400 24996 64424 24998
rect 64480 24996 64504 24998
rect 64560 24996 64584 24998
rect 64640 24996 64646 24998
rect 64338 24987 64646 24996
rect 64892 24750 64920 28727
rect 64984 28490 65012 28886
rect 65076 28762 65104 29718
rect 65064 28756 65116 28762
rect 65064 28698 65116 28704
rect 65168 28694 65196 31470
rect 65258 31036 65566 31045
rect 65258 31034 65264 31036
rect 65320 31034 65344 31036
rect 65400 31034 65424 31036
rect 65480 31034 65504 31036
rect 65560 31034 65566 31036
rect 65320 30982 65322 31034
rect 65502 30982 65504 31034
rect 65258 30980 65264 30982
rect 65320 30980 65344 30982
rect 65400 30980 65424 30982
rect 65480 30980 65504 30982
rect 65560 30980 65566 30982
rect 65258 30971 65566 30980
rect 65628 30258 65656 32166
rect 65812 31278 65840 34886
rect 65904 32434 65932 35634
rect 65996 33590 66024 35822
rect 66088 35698 66116 41006
rect 66444 37800 66496 37806
rect 66444 37742 66496 37748
rect 66260 36644 66312 36650
rect 66260 36586 66312 36592
rect 66272 35894 66300 36586
rect 66456 35894 66484 37742
rect 66534 36680 66590 36689
rect 66534 36615 66590 36624
rect 66180 35866 66300 35894
rect 66364 35866 66484 35894
rect 66076 35692 66128 35698
rect 66076 35634 66128 35640
rect 66076 35080 66128 35086
rect 66076 35022 66128 35028
rect 65984 33584 66036 33590
rect 65984 33526 66036 33532
rect 65984 33448 66036 33454
rect 65984 33390 66036 33396
rect 65996 32774 66024 33390
rect 66088 33046 66116 35022
rect 66076 33040 66128 33046
rect 66076 32982 66128 32988
rect 65984 32768 66036 32774
rect 65984 32710 66036 32716
rect 65984 32496 66036 32502
rect 65984 32438 66036 32444
rect 65892 32428 65944 32434
rect 65892 32370 65944 32376
rect 65996 31346 66024 32438
rect 66088 31346 66116 32982
rect 65984 31340 66036 31346
rect 65984 31282 66036 31288
rect 66076 31340 66128 31346
rect 66076 31282 66128 31288
rect 65800 31272 65852 31278
rect 66180 31226 66208 35866
rect 66260 33584 66312 33590
rect 66260 33526 66312 33532
rect 66272 32502 66300 33526
rect 66260 32496 66312 32502
rect 66260 32438 66312 32444
rect 65800 31214 65852 31220
rect 65708 31204 65760 31210
rect 65708 31146 65760 31152
rect 65904 31198 66208 31226
rect 65616 30252 65668 30258
rect 65616 30194 65668 30200
rect 65258 29948 65566 29957
rect 65258 29946 65264 29948
rect 65320 29946 65344 29948
rect 65400 29946 65424 29948
rect 65480 29946 65504 29948
rect 65560 29946 65566 29948
rect 65320 29894 65322 29946
rect 65502 29894 65504 29946
rect 65258 29892 65264 29894
rect 65320 29892 65344 29894
rect 65400 29892 65424 29894
rect 65480 29892 65504 29894
rect 65560 29892 65566 29894
rect 65258 29883 65566 29892
rect 65628 29646 65656 30194
rect 65720 29646 65748 31146
rect 65800 31136 65852 31142
rect 65800 31078 65852 31084
rect 65812 30870 65840 31078
rect 65800 30864 65852 30870
rect 65800 30806 65852 30812
rect 65616 29640 65668 29646
rect 65616 29582 65668 29588
rect 65708 29640 65760 29646
rect 65708 29582 65760 29588
rect 65258 28860 65566 28869
rect 65258 28858 65264 28860
rect 65320 28858 65344 28860
rect 65400 28858 65424 28860
rect 65480 28858 65504 28860
rect 65560 28858 65566 28860
rect 65320 28806 65322 28858
rect 65502 28806 65504 28858
rect 65258 28804 65264 28806
rect 65320 28804 65344 28806
rect 65400 28804 65424 28806
rect 65480 28804 65504 28806
rect 65560 28804 65566 28806
rect 65258 28795 65566 28804
rect 65156 28688 65208 28694
rect 65156 28630 65208 28636
rect 64972 28484 65024 28490
rect 64972 28426 65024 28432
rect 64984 26994 65012 28426
rect 65258 27772 65566 27781
rect 65258 27770 65264 27772
rect 65320 27770 65344 27772
rect 65400 27770 65424 27772
rect 65480 27770 65504 27772
rect 65560 27770 65566 27772
rect 65320 27718 65322 27770
rect 65502 27718 65504 27770
rect 65258 27716 65264 27718
rect 65320 27716 65344 27718
rect 65400 27716 65424 27718
rect 65480 27716 65504 27718
rect 65560 27716 65566 27718
rect 65258 27707 65566 27716
rect 65064 27056 65116 27062
rect 65064 26998 65116 27004
rect 64972 26988 65024 26994
rect 64972 26930 65024 26936
rect 64984 26586 65012 26930
rect 64972 26580 65024 26586
rect 64972 26522 65024 26528
rect 64972 26376 65024 26382
rect 64972 26318 65024 26324
rect 64880 24744 64932 24750
rect 64880 24686 64932 24692
rect 64984 24342 65012 26318
rect 65076 25906 65104 26998
rect 65628 26738 65656 29582
rect 65720 29170 65748 29582
rect 65708 29164 65760 29170
rect 65708 29106 65760 29112
rect 65720 26926 65748 29106
rect 65812 29034 65840 30806
rect 65800 29028 65852 29034
rect 65800 28970 65852 28976
rect 65708 26920 65760 26926
rect 65708 26862 65760 26868
rect 65800 26852 65852 26858
rect 65800 26794 65852 26800
rect 65628 26710 65748 26738
rect 65258 26684 65566 26693
rect 65258 26682 65264 26684
rect 65320 26682 65344 26684
rect 65400 26682 65424 26684
rect 65480 26682 65504 26684
rect 65560 26682 65566 26684
rect 65320 26630 65322 26682
rect 65502 26630 65504 26682
rect 65258 26628 65264 26630
rect 65320 26628 65344 26630
rect 65400 26628 65424 26630
rect 65480 26628 65504 26630
rect 65560 26628 65566 26630
rect 65258 26619 65566 26628
rect 65616 26580 65668 26586
rect 65616 26522 65668 26528
rect 65064 25900 65116 25906
rect 65064 25842 65116 25848
rect 65156 25900 65208 25906
rect 65156 25842 65208 25848
rect 65168 25294 65196 25842
rect 65258 25596 65566 25605
rect 65258 25594 65264 25596
rect 65320 25594 65344 25596
rect 65400 25594 65424 25596
rect 65480 25594 65504 25596
rect 65560 25594 65566 25596
rect 65320 25542 65322 25594
rect 65502 25542 65504 25594
rect 65258 25540 65264 25542
rect 65320 25540 65344 25542
rect 65400 25540 65424 25542
rect 65480 25540 65504 25542
rect 65560 25540 65566 25542
rect 65258 25531 65566 25540
rect 65064 25288 65116 25294
rect 65064 25230 65116 25236
rect 65156 25288 65208 25294
rect 65156 25230 65208 25236
rect 64236 24336 64288 24342
rect 64236 24278 64288 24284
rect 64972 24336 65024 24342
rect 64972 24278 65024 24284
rect 64338 23964 64646 23973
rect 64338 23962 64344 23964
rect 64400 23962 64424 23964
rect 64480 23962 64504 23964
rect 64560 23962 64584 23964
rect 64640 23962 64646 23964
rect 64400 23910 64402 23962
rect 64582 23910 64584 23962
rect 64338 23908 64344 23910
rect 64400 23908 64424 23910
rect 64480 23908 64504 23910
rect 64560 23908 64584 23910
rect 64640 23908 64646 23910
rect 64338 23899 64646 23908
rect 65076 23322 65104 25230
rect 65258 24508 65566 24517
rect 65258 24506 65264 24508
rect 65320 24506 65344 24508
rect 65400 24506 65424 24508
rect 65480 24506 65504 24508
rect 65560 24506 65566 24508
rect 65320 24454 65322 24506
rect 65502 24454 65504 24506
rect 65258 24452 65264 24454
rect 65320 24452 65344 24454
rect 65400 24452 65424 24454
rect 65480 24452 65504 24454
rect 65560 24452 65566 24454
rect 65258 24443 65566 24452
rect 65258 23420 65566 23429
rect 65258 23418 65264 23420
rect 65320 23418 65344 23420
rect 65400 23418 65424 23420
rect 65480 23418 65504 23420
rect 65560 23418 65566 23420
rect 65320 23366 65322 23418
rect 65502 23366 65504 23418
rect 65258 23364 65264 23366
rect 65320 23364 65344 23366
rect 65400 23364 65424 23366
rect 65480 23364 65504 23366
rect 65560 23364 65566 23366
rect 65258 23355 65566 23364
rect 65064 23316 65116 23322
rect 65064 23258 65116 23264
rect 64972 23180 65024 23186
rect 64972 23122 65024 23128
rect 64880 23044 64932 23050
rect 64880 22986 64932 22992
rect 64338 22876 64646 22885
rect 64338 22874 64344 22876
rect 64400 22874 64424 22876
rect 64480 22874 64504 22876
rect 64560 22874 64584 22876
rect 64640 22874 64646 22876
rect 64400 22822 64402 22874
rect 64582 22822 64584 22874
rect 64338 22820 64344 22822
rect 64400 22820 64424 22822
rect 64480 22820 64504 22822
rect 64560 22820 64584 22822
rect 64640 22820 64646 22822
rect 64338 22811 64646 22820
rect 64696 22024 64748 22030
rect 64696 21966 64748 21972
rect 64338 21788 64646 21797
rect 64338 21786 64344 21788
rect 64400 21786 64424 21788
rect 64480 21786 64504 21788
rect 64560 21786 64584 21788
rect 64640 21786 64646 21788
rect 64400 21734 64402 21786
rect 64582 21734 64584 21786
rect 64338 21732 64344 21734
rect 64400 21732 64424 21734
rect 64480 21732 64504 21734
rect 64560 21732 64584 21734
rect 64640 21732 64646 21734
rect 64338 21723 64646 21732
rect 64708 21146 64736 21966
rect 64696 21140 64748 21146
rect 64696 21082 64748 21088
rect 64156 20726 64276 20754
rect 64144 20596 64196 20602
rect 64144 20538 64196 20544
rect 64052 19916 64104 19922
rect 64052 19858 64104 19864
rect 64064 18290 64092 19858
rect 64052 18284 64104 18290
rect 64052 18226 64104 18232
rect 63880 16546 64000 16574
rect 63880 14958 63908 16546
rect 63868 14952 63920 14958
rect 63868 14894 63920 14900
rect 63880 13326 63908 14894
rect 63868 13320 63920 13326
rect 63868 13262 63920 13268
rect 63880 12238 63908 13262
rect 63868 12232 63920 12238
rect 63868 12174 63920 12180
rect 63880 8974 63908 12174
rect 63960 11552 64012 11558
rect 63960 11494 64012 11500
rect 63868 8968 63920 8974
rect 63868 8910 63920 8916
rect 63776 6860 63828 6866
rect 63776 6802 63828 6808
rect 63788 3398 63816 6802
rect 63880 5234 63908 8910
rect 63972 6390 64000 11494
rect 64064 7954 64092 18226
rect 64156 15366 64184 20538
rect 64248 17882 64276 20726
rect 64338 20700 64646 20709
rect 64338 20698 64344 20700
rect 64400 20698 64424 20700
rect 64480 20698 64504 20700
rect 64560 20698 64584 20700
rect 64640 20698 64646 20700
rect 64400 20646 64402 20698
rect 64582 20646 64584 20698
rect 64338 20644 64344 20646
rect 64400 20644 64424 20646
rect 64480 20644 64504 20646
rect 64560 20644 64584 20646
rect 64640 20644 64646 20646
rect 64338 20635 64646 20644
rect 64696 19848 64748 19854
rect 64696 19790 64748 19796
rect 64338 19612 64646 19621
rect 64338 19610 64344 19612
rect 64400 19610 64424 19612
rect 64480 19610 64504 19612
rect 64560 19610 64584 19612
rect 64640 19610 64646 19612
rect 64400 19558 64402 19610
rect 64582 19558 64584 19610
rect 64338 19556 64344 19558
rect 64400 19556 64424 19558
rect 64480 19556 64504 19558
rect 64560 19556 64584 19558
rect 64640 19556 64646 19558
rect 64338 19547 64646 19556
rect 64708 19514 64736 19790
rect 64696 19508 64748 19514
rect 64696 19450 64748 19456
rect 64892 19334 64920 22986
rect 64984 22778 65012 23122
rect 65628 23118 65656 26522
rect 65720 25906 65748 26710
rect 65708 25900 65760 25906
rect 65708 25842 65760 25848
rect 65812 25294 65840 26794
rect 65800 25288 65852 25294
rect 65800 25230 65852 25236
rect 65812 24070 65840 25230
rect 65800 24064 65852 24070
rect 65800 24006 65852 24012
rect 65616 23112 65668 23118
rect 65616 23054 65668 23060
rect 64972 22772 65024 22778
rect 64972 22714 65024 22720
rect 65258 22332 65566 22341
rect 65258 22330 65264 22332
rect 65320 22330 65344 22332
rect 65400 22330 65424 22332
rect 65480 22330 65504 22332
rect 65560 22330 65566 22332
rect 65320 22278 65322 22330
rect 65502 22278 65504 22330
rect 65258 22276 65264 22278
rect 65320 22276 65344 22278
rect 65400 22276 65424 22278
rect 65480 22276 65504 22278
rect 65560 22276 65566 22278
rect 65258 22267 65566 22276
rect 65616 21412 65668 21418
rect 65616 21354 65668 21360
rect 64972 21344 65024 21350
rect 64972 21286 65024 21292
rect 64984 21146 65012 21286
rect 65258 21244 65566 21253
rect 65258 21242 65264 21244
rect 65320 21242 65344 21244
rect 65400 21242 65424 21244
rect 65480 21242 65504 21244
rect 65560 21242 65566 21244
rect 65320 21190 65322 21242
rect 65502 21190 65504 21242
rect 65258 21188 65264 21190
rect 65320 21188 65344 21190
rect 65400 21188 65424 21190
rect 65480 21188 65504 21190
rect 65560 21188 65566 21190
rect 65258 21179 65566 21188
rect 64972 21140 65024 21146
rect 64972 21082 65024 21088
rect 65156 21072 65208 21078
rect 65156 21014 65208 21020
rect 65064 20528 65116 20534
rect 65064 20470 65116 20476
rect 64972 20256 65024 20262
rect 64972 20198 65024 20204
rect 64800 19306 64920 19334
rect 64696 18624 64748 18630
rect 64696 18566 64748 18572
rect 64338 18524 64646 18533
rect 64338 18522 64344 18524
rect 64400 18522 64424 18524
rect 64480 18522 64504 18524
rect 64560 18522 64584 18524
rect 64640 18522 64646 18524
rect 64400 18470 64402 18522
rect 64582 18470 64584 18522
rect 64338 18468 64344 18470
rect 64400 18468 64424 18470
rect 64480 18468 64504 18470
rect 64560 18468 64584 18470
rect 64640 18468 64646 18470
rect 64338 18459 64646 18468
rect 64708 18290 64736 18566
rect 64696 18284 64748 18290
rect 64696 18226 64748 18232
rect 64236 17876 64288 17882
rect 64236 17818 64288 17824
rect 64248 17338 64276 17818
rect 64338 17436 64646 17445
rect 64338 17434 64344 17436
rect 64400 17434 64424 17436
rect 64480 17434 64504 17436
rect 64560 17434 64584 17436
rect 64640 17434 64646 17436
rect 64400 17382 64402 17434
rect 64582 17382 64584 17434
rect 64338 17380 64344 17382
rect 64400 17380 64424 17382
rect 64480 17380 64504 17382
rect 64560 17380 64584 17382
rect 64640 17380 64646 17382
rect 64338 17371 64646 17380
rect 64236 17332 64288 17338
rect 64236 17274 64288 17280
rect 64800 16574 64828 19306
rect 64880 17672 64932 17678
rect 64880 17614 64932 17620
rect 64708 16546 64828 16574
rect 64338 16348 64646 16357
rect 64338 16346 64344 16348
rect 64400 16346 64424 16348
rect 64480 16346 64504 16348
rect 64560 16346 64584 16348
rect 64640 16346 64646 16348
rect 64400 16294 64402 16346
rect 64582 16294 64584 16346
rect 64338 16292 64344 16294
rect 64400 16292 64424 16294
rect 64480 16292 64504 16294
rect 64560 16292 64584 16294
rect 64640 16292 64646 16294
rect 64338 16283 64646 16292
rect 64708 16232 64736 16546
rect 64892 16250 64920 17614
rect 64984 16794 65012 20198
rect 65076 19310 65104 20470
rect 65064 19304 65116 19310
rect 65064 19246 65116 19252
rect 65064 18760 65116 18766
rect 65064 18702 65116 18708
rect 65076 17882 65104 18702
rect 65064 17876 65116 17882
rect 65064 17818 65116 17824
rect 65168 17610 65196 21014
rect 65628 20942 65656 21354
rect 65616 20936 65668 20942
rect 65616 20878 65668 20884
rect 65258 20156 65566 20165
rect 65258 20154 65264 20156
rect 65320 20154 65344 20156
rect 65400 20154 65424 20156
rect 65480 20154 65504 20156
rect 65560 20154 65566 20156
rect 65320 20102 65322 20154
rect 65502 20102 65504 20154
rect 65258 20100 65264 20102
rect 65320 20100 65344 20102
rect 65400 20100 65424 20102
rect 65480 20100 65504 20102
rect 65560 20100 65566 20102
rect 65258 20091 65566 20100
rect 65628 19378 65656 20878
rect 65708 20460 65760 20466
rect 65708 20402 65760 20408
rect 65616 19372 65668 19378
rect 65616 19314 65668 19320
rect 65258 19068 65566 19077
rect 65258 19066 65264 19068
rect 65320 19066 65344 19068
rect 65400 19066 65424 19068
rect 65480 19066 65504 19068
rect 65560 19066 65566 19068
rect 65320 19014 65322 19066
rect 65502 19014 65504 19066
rect 65258 19012 65264 19014
rect 65320 19012 65344 19014
rect 65400 19012 65424 19014
rect 65480 19012 65504 19014
rect 65560 19012 65566 19014
rect 65258 19003 65566 19012
rect 65628 18766 65656 19314
rect 65616 18760 65668 18766
rect 65616 18702 65668 18708
rect 65258 17980 65566 17989
rect 65258 17978 65264 17980
rect 65320 17978 65344 17980
rect 65400 17978 65424 17980
rect 65480 17978 65504 17980
rect 65560 17978 65566 17980
rect 65320 17926 65322 17978
rect 65502 17926 65504 17978
rect 65258 17924 65264 17926
rect 65320 17924 65344 17926
rect 65400 17924 65424 17926
rect 65480 17924 65504 17926
rect 65560 17924 65566 17926
rect 65258 17915 65566 17924
rect 65156 17604 65208 17610
rect 65156 17546 65208 17552
rect 65258 16892 65566 16901
rect 65258 16890 65264 16892
rect 65320 16890 65344 16892
rect 65400 16890 65424 16892
rect 65480 16890 65504 16892
rect 65560 16890 65566 16892
rect 65320 16838 65322 16890
rect 65502 16838 65504 16890
rect 65258 16836 65264 16838
rect 65320 16836 65344 16838
rect 65400 16836 65424 16838
rect 65480 16836 65504 16838
rect 65560 16836 65566 16838
rect 65258 16827 65566 16836
rect 64972 16788 65024 16794
rect 64972 16730 65024 16736
rect 65156 16720 65208 16726
rect 64970 16688 65026 16697
rect 64970 16623 65026 16632
rect 65076 16668 65156 16674
rect 65076 16662 65208 16668
rect 65076 16646 65196 16662
rect 64616 16204 64736 16232
rect 64880 16244 64932 16250
rect 64616 16046 64644 16204
rect 64880 16186 64932 16192
rect 64788 16176 64840 16182
rect 64788 16118 64840 16124
rect 64604 16040 64656 16046
rect 64604 15982 64656 15988
rect 64616 15706 64644 15982
rect 64604 15700 64656 15706
rect 64604 15642 64656 15648
rect 64144 15360 64196 15366
rect 64144 15302 64196 15308
rect 64338 15260 64646 15269
rect 64338 15258 64344 15260
rect 64400 15258 64424 15260
rect 64480 15258 64504 15260
rect 64560 15258 64584 15260
rect 64640 15258 64646 15260
rect 64400 15206 64402 15258
rect 64582 15206 64584 15258
rect 64338 15204 64344 15206
rect 64400 15204 64424 15206
rect 64480 15204 64504 15206
rect 64560 15204 64584 15206
rect 64640 15204 64646 15206
rect 64142 15192 64198 15201
rect 64338 15195 64646 15204
rect 64142 15127 64198 15136
rect 64052 7948 64104 7954
rect 64052 7890 64104 7896
rect 63960 6384 64012 6390
rect 63960 6326 64012 6332
rect 63960 5704 64012 5710
rect 63960 5646 64012 5652
rect 63868 5228 63920 5234
rect 63868 5170 63920 5176
rect 63972 3534 64000 5646
rect 64064 4690 64092 7890
rect 64156 7546 64184 15127
rect 64800 15026 64828 16118
rect 64788 15020 64840 15026
rect 64788 14962 64840 14968
rect 64338 14172 64646 14181
rect 64338 14170 64344 14172
rect 64400 14170 64424 14172
rect 64480 14170 64504 14172
rect 64560 14170 64584 14172
rect 64640 14170 64646 14172
rect 64400 14118 64402 14170
rect 64582 14118 64584 14170
rect 64338 14116 64344 14118
rect 64400 14116 64424 14118
rect 64480 14116 64504 14118
rect 64560 14116 64584 14118
rect 64640 14116 64646 14118
rect 64338 14107 64646 14116
rect 64236 13456 64288 13462
rect 64236 13398 64288 13404
rect 64248 11898 64276 13398
rect 64338 13084 64646 13093
rect 64338 13082 64344 13084
rect 64400 13082 64424 13084
rect 64480 13082 64504 13084
rect 64560 13082 64584 13084
rect 64640 13082 64646 13084
rect 64400 13030 64402 13082
rect 64582 13030 64584 13082
rect 64338 13028 64344 13030
rect 64400 13028 64424 13030
rect 64480 13028 64504 13030
rect 64560 13028 64584 13030
rect 64640 13028 64646 13030
rect 64338 13019 64646 13028
rect 64696 12232 64748 12238
rect 64696 12174 64748 12180
rect 64338 11996 64646 12005
rect 64338 11994 64344 11996
rect 64400 11994 64424 11996
rect 64480 11994 64504 11996
rect 64560 11994 64584 11996
rect 64640 11994 64646 11996
rect 64400 11942 64402 11994
rect 64582 11942 64584 11994
rect 64338 11940 64344 11942
rect 64400 11940 64424 11942
rect 64480 11940 64504 11942
rect 64560 11940 64584 11942
rect 64640 11940 64646 11942
rect 64338 11931 64646 11940
rect 64236 11892 64288 11898
rect 64236 11834 64288 11840
rect 64708 11354 64736 12174
rect 64696 11348 64748 11354
rect 64696 11290 64748 11296
rect 64338 10908 64646 10917
rect 64338 10906 64344 10908
rect 64400 10906 64424 10908
rect 64480 10906 64504 10908
rect 64560 10906 64584 10908
rect 64640 10906 64646 10908
rect 64400 10854 64402 10906
rect 64582 10854 64584 10906
rect 64338 10852 64344 10854
rect 64400 10852 64424 10854
rect 64480 10852 64504 10854
rect 64560 10852 64584 10854
rect 64640 10852 64646 10854
rect 64338 10843 64646 10852
rect 64892 10674 64920 16186
rect 64984 15178 65012 16623
rect 65076 16574 65104 16646
rect 65076 16546 65196 16574
rect 64984 15150 65104 15178
rect 65076 14890 65104 15150
rect 65064 14884 65116 14890
rect 65064 14826 65116 14832
rect 64972 12640 65024 12646
rect 64972 12582 65024 12588
rect 64984 11694 65012 12582
rect 64972 11688 65024 11694
rect 64972 11630 65024 11636
rect 64880 10668 64932 10674
rect 64880 10610 64932 10616
rect 64892 10554 64920 10610
rect 64892 10526 65012 10554
rect 64788 10464 64840 10470
rect 64788 10406 64840 10412
rect 64880 10464 64932 10470
rect 64880 10406 64932 10412
rect 64338 9820 64646 9829
rect 64338 9818 64344 9820
rect 64400 9818 64424 9820
rect 64480 9818 64504 9820
rect 64560 9818 64584 9820
rect 64640 9818 64646 9820
rect 64400 9766 64402 9818
rect 64582 9766 64584 9818
rect 64338 9764 64344 9766
rect 64400 9764 64424 9766
rect 64480 9764 64504 9766
rect 64560 9764 64584 9766
rect 64640 9764 64646 9766
rect 64338 9755 64646 9764
rect 64696 8968 64748 8974
rect 64696 8910 64748 8916
rect 64338 8732 64646 8741
rect 64338 8730 64344 8732
rect 64400 8730 64424 8732
rect 64480 8730 64504 8732
rect 64560 8730 64584 8732
rect 64640 8730 64646 8732
rect 64400 8678 64402 8730
rect 64582 8678 64584 8730
rect 64338 8676 64344 8678
rect 64400 8676 64424 8678
rect 64480 8676 64504 8678
rect 64560 8676 64584 8678
rect 64640 8676 64646 8678
rect 64338 8667 64646 8676
rect 64708 8634 64736 8910
rect 64696 8628 64748 8634
rect 64696 8570 64748 8576
rect 64696 7880 64748 7886
rect 64696 7822 64748 7828
rect 64338 7644 64646 7653
rect 64338 7642 64344 7644
rect 64400 7642 64424 7644
rect 64480 7642 64504 7644
rect 64560 7642 64584 7644
rect 64640 7642 64646 7644
rect 64400 7590 64402 7642
rect 64582 7590 64584 7642
rect 64338 7588 64344 7590
rect 64400 7588 64424 7590
rect 64480 7588 64504 7590
rect 64560 7588 64584 7590
rect 64640 7588 64646 7590
rect 64338 7579 64646 7588
rect 64708 7546 64736 7822
rect 64144 7540 64196 7546
rect 64144 7482 64196 7488
rect 64696 7540 64748 7546
rect 64696 7482 64748 7488
rect 64156 7002 64184 7482
rect 64800 7410 64828 10406
rect 64892 10062 64920 10406
rect 64984 10130 65012 10526
rect 64972 10124 65024 10130
rect 64972 10066 65024 10072
rect 64880 10056 64932 10062
rect 64880 9998 64932 10004
rect 64984 9466 65012 10066
rect 64892 9438 65012 9466
rect 64788 7404 64840 7410
rect 64788 7346 64840 7352
rect 64144 6996 64196 7002
rect 64144 6938 64196 6944
rect 64156 6458 64184 6938
rect 64892 6798 64920 9438
rect 64972 9376 65024 9382
rect 64972 9318 65024 9324
rect 64984 7342 65012 9318
rect 65076 8514 65104 14826
rect 65168 14822 65196 16546
rect 65258 15804 65566 15813
rect 65258 15802 65264 15804
rect 65320 15802 65344 15804
rect 65400 15802 65424 15804
rect 65480 15802 65504 15804
rect 65560 15802 65566 15804
rect 65320 15750 65322 15802
rect 65502 15750 65504 15802
rect 65258 15748 65264 15750
rect 65320 15748 65344 15750
rect 65400 15748 65424 15750
rect 65480 15748 65504 15750
rect 65560 15748 65566 15750
rect 65258 15739 65566 15748
rect 65156 14816 65208 14822
rect 65156 14758 65208 14764
rect 65258 14716 65566 14725
rect 65258 14714 65264 14716
rect 65320 14714 65344 14716
rect 65400 14714 65424 14716
rect 65480 14714 65504 14716
rect 65560 14714 65566 14716
rect 65320 14662 65322 14714
rect 65502 14662 65504 14714
rect 65258 14660 65264 14662
rect 65320 14660 65344 14662
rect 65400 14660 65424 14662
rect 65480 14660 65504 14662
rect 65560 14660 65566 14662
rect 65258 14651 65566 14660
rect 65628 13818 65656 18702
rect 65720 17746 65748 20402
rect 65812 20398 65840 24006
rect 65904 20602 65932 31198
rect 66364 31090 66392 35866
rect 66444 33380 66496 33386
rect 66444 33322 66496 33328
rect 66088 31062 66392 31090
rect 65984 30592 66036 30598
rect 65984 30534 66036 30540
rect 65996 30190 66024 30534
rect 65984 30184 66036 30190
rect 65984 30126 66036 30132
rect 65996 28626 66024 30126
rect 65984 28620 66036 28626
rect 65984 28562 66036 28568
rect 65984 26240 66036 26246
rect 65984 26182 66036 26188
rect 65996 25838 66024 26182
rect 65984 25832 66036 25838
rect 65984 25774 66036 25780
rect 65996 23254 66024 25774
rect 65984 23248 66036 23254
rect 65984 23190 66036 23196
rect 66088 21078 66116 31062
rect 66168 29028 66220 29034
rect 66168 28970 66220 28976
rect 66180 26518 66208 28970
rect 66168 26512 66220 26518
rect 66168 26454 66220 26460
rect 66456 26234 66484 33322
rect 66364 26206 66484 26234
rect 66364 22234 66392 26206
rect 66548 23186 66576 36615
rect 66536 23180 66588 23186
rect 66536 23122 66588 23128
rect 66352 22228 66404 22234
rect 66352 22170 66404 22176
rect 66168 22160 66220 22166
rect 66168 22102 66220 22108
rect 66076 21072 66128 21078
rect 66076 21014 66128 21020
rect 65892 20596 65944 20602
rect 65892 20538 65944 20544
rect 65800 20392 65852 20398
rect 65800 20334 65852 20340
rect 65984 19712 66036 19718
rect 65984 19654 66036 19660
rect 65996 19310 66024 19654
rect 65984 19304 66036 19310
rect 65984 19246 66036 19252
rect 65800 18760 65852 18766
rect 65800 18702 65852 18708
rect 65812 18086 65840 18702
rect 65800 18080 65852 18086
rect 65800 18022 65852 18028
rect 65812 17814 65840 18022
rect 65800 17808 65852 17814
rect 65800 17750 65852 17756
rect 65708 17740 65760 17746
rect 65708 17682 65760 17688
rect 65708 17604 65760 17610
rect 65708 17546 65760 17552
rect 65168 13790 65656 13818
rect 65168 11762 65196 13790
rect 65258 13628 65566 13637
rect 65258 13626 65264 13628
rect 65320 13626 65344 13628
rect 65400 13626 65424 13628
rect 65480 13626 65504 13628
rect 65560 13626 65566 13628
rect 65320 13574 65322 13626
rect 65502 13574 65504 13626
rect 65258 13572 65264 13574
rect 65320 13572 65344 13574
rect 65400 13572 65424 13574
rect 65480 13572 65504 13574
rect 65560 13572 65566 13574
rect 65258 13563 65566 13572
rect 65720 13530 65748 17546
rect 65892 16448 65944 16454
rect 65892 16390 65944 16396
rect 65904 16114 65932 16390
rect 65996 16182 66024 19246
rect 66088 16697 66116 21014
rect 66180 20806 66208 22102
rect 66364 21554 66392 22170
rect 66352 21548 66404 21554
rect 66352 21490 66404 21496
rect 66168 20800 66220 20806
rect 66168 20742 66220 20748
rect 66180 19990 66208 20742
rect 66168 19984 66220 19990
rect 66168 19926 66220 19932
rect 66180 18154 66208 19926
rect 66168 18148 66220 18154
rect 66168 18090 66220 18096
rect 66074 16688 66130 16697
rect 66074 16623 66130 16632
rect 66076 16448 66128 16454
rect 66076 16390 66128 16396
rect 65984 16176 66036 16182
rect 65984 16118 66036 16124
rect 65892 16108 65944 16114
rect 65892 16050 65944 16056
rect 66088 16046 66116 16390
rect 66076 16040 66128 16046
rect 66076 15982 66128 15988
rect 65800 14816 65852 14822
rect 65800 14758 65852 14764
rect 65708 13524 65760 13530
rect 65708 13466 65760 13472
rect 65616 13456 65668 13462
rect 65616 13398 65668 13404
rect 65258 12540 65566 12549
rect 65258 12538 65264 12540
rect 65320 12538 65344 12540
rect 65400 12538 65424 12540
rect 65480 12538 65504 12540
rect 65560 12538 65566 12540
rect 65320 12486 65322 12538
rect 65502 12486 65504 12538
rect 65258 12484 65264 12486
rect 65320 12484 65344 12486
rect 65400 12484 65424 12486
rect 65480 12484 65504 12486
rect 65560 12484 65566 12486
rect 65258 12475 65566 12484
rect 65628 12374 65656 13398
rect 65720 12850 65748 13466
rect 65708 12844 65760 12850
rect 65708 12786 65760 12792
rect 65616 12368 65668 12374
rect 65616 12310 65668 12316
rect 65156 11756 65208 11762
rect 65156 11698 65208 11704
rect 65168 11150 65196 11698
rect 65258 11452 65566 11461
rect 65258 11450 65264 11452
rect 65320 11450 65344 11452
rect 65400 11450 65424 11452
rect 65480 11450 65504 11452
rect 65560 11450 65566 11452
rect 65320 11398 65322 11450
rect 65502 11398 65504 11450
rect 65258 11396 65264 11398
rect 65320 11396 65344 11398
rect 65400 11396 65424 11398
rect 65480 11396 65504 11398
rect 65560 11396 65566 11398
rect 65258 11387 65566 11396
rect 65156 11144 65208 11150
rect 65156 11086 65208 11092
rect 65168 8650 65196 11086
rect 65258 10364 65566 10373
rect 65258 10362 65264 10364
rect 65320 10362 65344 10364
rect 65400 10362 65424 10364
rect 65480 10362 65504 10364
rect 65560 10362 65566 10364
rect 65320 10310 65322 10362
rect 65502 10310 65504 10362
rect 65258 10308 65264 10310
rect 65320 10308 65344 10310
rect 65400 10308 65424 10310
rect 65480 10308 65504 10310
rect 65560 10308 65566 10310
rect 65258 10299 65566 10308
rect 65258 9276 65566 9285
rect 65258 9274 65264 9276
rect 65320 9274 65344 9276
rect 65400 9274 65424 9276
rect 65480 9274 65504 9276
rect 65560 9274 65566 9276
rect 65320 9222 65322 9274
rect 65502 9222 65504 9274
rect 65258 9220 65264 9222
rect 65320 9220 65344 9222
rect 65400 9220 65424 9222
rect 65480 9220 65504 9222
rect 65560 9220 65566 9222
rect 65258 9211 65566 9220
rect 65628 9110 65656 12310
rect 65720 10266 65748 12786
rect 65812 10606 65840 14758
rect 66180 13462 66208 18090
rect 66364 17882 66392 21490
rect 66352 17876 66404 17882
rect 66352 17818 66404 17824
rect 66444 16108 66496 16114
rect 66444 16050 66496 16056
rect 66168 13456 66220 13462
rect 66168 13398 66220 13404
rect 66352 12232 66404 12238
rect 66352 12174 66404 12180
rect 66364 11286 66392 12174
rect 66352 11280 66404 11286
rect 66352 11222 66404 11228
rect 66168 11212 66220 11218
rect 66168 11154 66220 11160
rect 65800 10600 65852 10606
rect 65800 10542 65852 10548
rect 65708 10260 65760 10266
rect 65708 10202 65760 10208
rect 65984 10056 66036 10062
rect 65984 9998 66036 10004
rect 65708 9920 65760 9926
rect 65708 9862 65760 9868
rect 65616 9104 65668 9110
rect 65616 9046 65668 9052
rect 65168 8622 65288 8650
rect 65076 8486 65196 8514
rect 65260 8498 65288 8622
rect 65064 8424 65116 8430
rect 65064 8366 65116 8372
rect 64972 7336 65024 7342
rect 64972 7278 65024 7284
rect 64880 6792 64932 6798
rect 64880 6734 64932 6740
rect 64236 6656 64288 6662
rect 64236 6598 64288 6604
rect 64144 6452 64196 6458
rect 64144 6394 64196 6400
rect 64142 5944 64198 5953
rect 64142 5879 64144 5888
rect 64196 5879 64198 5888
rect 64144 5850 64196 5856
rect 64248 4758 64276 6598
rect 64338 6556 64646 6565
rect 64338 6554 64344 6556
rect 64400 6554 64424 6556
rect 64480 6554 64504 6556
rect 64560 6554 64584 6556
rect 64640 6554 64646 6556
rect 64400 6502 64402 6554
rect 64582 6502 64584 6554
rect 64338 6500 64344 6502
rect 64400 6500 64424 6502
rect 64480 6500 64504 6502
rect 64560 6500 64584 6502
rect 64640 6500 64646 6502
rect 64338 6491 64646 6500
rect 64892 6322 64920 6734
rect 65076 6730 65104 8366
rect 65064 6724 65116 6730
rect 65064 6666 65116 6672
rect 64880 6316 64932 6322
rect 64880 6258 64932 6264
rect 64696 6112 64748 6118
rect 64694 6080 64696 6089
rect 64748 6080 64750 6089
rect 64892 6066 64920 6258
rect 64694 6015 64750 6024
rect 64800 6038 64920 6066
rect 64708 5914 64736 6015
rect 64696 5908 64748 5914
rect 64696 5850 64748 5856
rect 64800 5778 64828 6038
rect 64880 5908 64932 5914
rect 64880 5850 64932 5856
rect 64788 5772 64840 5778
rect 64788 5714 64840 5720
rect 64696 5704 64748 5710
rect 64696 5646 64748 5652
rect 64338 5468 64646 5477
rect 64338 5466 64344 5468
rect 64400 5466 64424 5468
rect 64480 5466 64504 5468
rect 64560 5466 64584 5468
rect 64640 5466 64646 5468
rect 64400 5414 64402 5466
rect 64582 5414 64584 5466
rect 64338 5412 64344 5414
rect 64400 5412 64424 5414
rect 64480 5412 64504 5414
rect 64560 5412 64584 5414
rect 64640 5412 64646 5414
rect 64338 5403 64646 5412
rect 64236 4752 64288 4758
rect 64236 4694 64288 4700
rect 64052 4684 64104 4690
rect 64052 4626 64104 4632
rect 64064 4010 64092 4626
rect 64338 4380 64646 4389
rect 64338 4378 64344 4380
rect 64400 4378 64424 4380
rect 64480 4378 64504 4380
rect 64560 4378 64584 4380
rect 64640 4378 64646 4380
rect 64400 4326 64402 4378
rect 64582 4326 64584 4378
rect 64338 4324 64344 4326
rect 64400 4324 64424 4326
rect 64480 4324 64504 4326
rect 64560 4324 64584 4326
rect 64640 4324 64646 4326
rect 64338 4315 64646 4324
rect 64236 4276 64288 4282
rect 64236 4218 64288 4224
rect 64052 4004 64104 4010
rect 64052 3946 64104 3952
rect 64144 4004 64196 4010
rect 64144 3946 64196 3952
rect 63960 3528 64012 3534
rect 63960 3470 64012 3476
rect 63776 3392 63828 3398
rect 63776 3334 63828 3340
rect 64064 3058 64092 3946
rect 64156 3738 64184 3946
rect 64144 3732 64196 3738
rect 64144 3674 64196 3680
rect 64248 3670 64276 4218
rect 64236 3664 64288 3670
rect 64236 3606 64288 3612
rect 64248 3210 64276 3606
rect 64708 3466 64736 5646
rect 64788 5568 64840 5574
rect 64788 5510 64840 5516
rect 64800 5234 64828 5510
rect 64788 5228 64840 5234
rect 64788 5170 64840 5176
rect 64696 3460 64748 3466
rect 64696 3402 64748 3408
rect 64788 3392 64840 3398
rect 64788 3334 64840 3340
rect 64338 3292 64646 3301
rect 64338 3290 64344 3292
rect 64400 3290 64424 3292
rect 64480 3290 64504 3292
rect 64560 3290 64584 3292
rect 64640 3290 64646 3292
rect 64400 3238 64402 3290
rect 64582 3238 64584 3290
rect 64338 3236 64344 3238
rect 64400 3236 64424 3238
rect 64480 3236 64504 3238
rect 64560 3236 64584 3238
rect 64640 3236 64646 3238
rect 64338 3227 64646 3236
rect 64156 3194 64276 3210
rect 64144 3188 64276 3194
rect 64196 3182 64276 3188
rect 64144 3130 64196 3136
rect 64052 3052 64104 3058
rect 64052 2994 64104 3000
rect 64328 2916 64380 2922
rect 64328 2858 64380 2864
rect 64340 2650 64368 2858
rect 64328 2644 64380 2650
rect 64328 2586 64380 2592
rect 64800 2446 64828 3334
rect 64788 2440 64840 2446
rect 64788 2382 64840 2388
rect 64892 2310 64920 5850
rect 65064 5772 65116 5778
rect 65064 5714 65116 5720
rect 64972 5636 65024 5642
rect 64972 5578 65024 5584
rect 64984 3534 65012 5578
rect 64972 3528 65024 3534
rect 64972 3470 65024 3476
rect 64972 2508 65024 2514
rect 64972 2450 65024 2456
rect 64880 2304 64932 2310
rect 64880 2246 64932 2252
rect 64338 2204 64646 2213
rect 64338 2202 64344 2204
rect 64400 2202 64424 2204
rect 64480 2202 64504 2204
rect 64560 2202 64584 2204
rect 64640 2202 64646 2204
rect 64400 2150 64402 2202
rect 64582 2150 64584 2202
rect 64338 2148 64344 2150
rect 64400 2148 64424 2150
rect 64480 2148 64504 2150
rect 64560 2148 64584 2150
rect 64640 2148 64646 2150
rect 64338 2139 64646 2148
rect 64694 2000 64750 2009
rect 64694 1935 64750 1944
rect 64708 1902 64736 1935
rect 64696 1896 64748 1902
rect 63040 1838 63092 1844
rect 63498 1864 63554 1873
rect 64696 1838 64748 1844
rect 63498 1799 63554 1808
rect 62854 1592 62910 1601
rect 62854 1527 62910 1536
rect 64708 1358 64736 1838
rect 64696 1352 64748 1358
rect 62578 1320 62634 1329
rect 64696 1294 64748 1300
rect 62578 1255 62634 1264
rect 64338 1116 64646 1125
rect 64338 1114 64344 1116
rect 64400 1114 64424 1116
rect 64480 1114 64504 1116
rect 64560 1114 64584 1116
rect 64640 1114 64646 1116
rect 64400 1062 64402 1114
rect 64582 1062 64584 1114
rect 64338 1060 64344 1062
rect 64400 1060 64424 1062
rect 64480 1060 64504 1062
rect 64560 1060 64584 1062
rect 64640 1060 64646 1062
rect 64338 1051 64646 1060
rect 64984 1018 65012 2450
rect 65076 2106 65104 5714
rect 65168 4010 65196 8486
rect 65248 8492 65300 8498
rect 65248 8434 65300 8440
rect 65258 8188 65566 8197
rect 65258 8186 65264 8188
rect 65320 8186 65344 8188
rect 65400 8186 65424 8188
rect 65480 8186 65504 8188
rect 65560 8186 65566 8188
rect 65320 8134 65322 8186
rect 65502 8134 65504 8186
rect 65258 8132 65264 8134
rect 65320 8132 65344 8134
rect 65400 8132 65424 8134
rect 65480 8132 65504 8134
rect 65560 8132 65566 8134
rect 65258 8123 65566 8132
rect 65628 8022 65656 9046
rect 65616 8016 65668 8022
rect 65616 7958 65668 7964
rect 65616 7200 65668 7206
rect 65616 7142 65668 7148
rect 65258 7100 65566 7109
rect 65258 7098 65264 7100
rect 65320 7098 65344 7100
rect 65400 7098 65424 7100
rect 65480 7098 65504 7100
rect 65560 7098 65566 7100
rect 65320 7046 65322 7098
rect 65502 7046 65504 7098
rect 65258 7044 65264 7046
rect 65320 7044 65344 7046
rect 65400 7044 65424 7046
rect 65480 7044 65504 7046
rect 65560 7044 65566 7046
rect 65258 7035 65566 7044
rect 65628 7002 65656 7142
rect 65616 6996 65668 7002
rect 65616 6938 65668 6944
rect 65720 6866 65748 9862
rect 65800 9512 65852 9518
rect 65800 9454 65852 9460
rect 65812 8090 65840 9454
rect 65996 8838 66024 9998
rect 65984 8832 66036 8838
rect 65984 8774 66036 8780
rect 65996 8498 66024 8774
rect 65892 8492 65944 8498
rect 65892 8434 65944 8440
rect 65984 8492 66036 8498
rect 65984 8434 66036 8440
rect 65800 8084 65852 8090
rect 65800 8026 65852 8032
rect 65812 6934 65840 8026
rect 65904 7410 65932 8434
rect 66076 8016 66128 8022
rect 66076 7958 66128 7964
rect 65892 7404 65944 7410
rect 65892 7346 65944 7352
rect 65800 6928 65852 6934
rect 65800 6870 65852 6876
rect 65708 6860 65760 6866
rect 65708 6802 65760 6808
rect 65800 6792 65852 6798
rect 65904 6746 65932 7346
rect 65984 7336 66036 7342
rect 65984 7278 66036 7284
rect 65852 6740 65932 6746
rect 65800 6734 65932 6740
rect 65812 6718 65932 6734
rect 65258 6012 65566 6021
rect 65258 6010 65264 6012
rect 65320 6010 65344 6012
rect 65400 6010 65424 6012
rect 65480 6010 65504 6012
rect 65560 6010 65566 6012
rect 65320 5958 65322 6010
rect 65502 5958 65504 6010
rect 65258 5956 65264 5958
rect 65320 5956 65344 5958
rect 65400 5956 65424 5958
rect 65480 5956 65504 5958
rect 65560 5956 65566 5958
rect 65258 5947 65566 5956
rect 65812 5914 65840 6718
rect 65996 6254 66024 7278
rect 65984 6248 66036 6254
rect 65984 6190 66036 6196
rect 65432 5908 65484 5914
rect 65432 5850 65484 5856
rect 65800 5908 65852 5914
rect 65800 5850 65852 5856
rect 65444 5710 65472 5850
rect 65708 5840 65760 5846
rect 65708 5782 65760 5788
rect 65432 5704 65484 5710
rect 65432 5646 65484 5652
rect 65616 5160 65668 5166
rect 65616 5102 65668 5108
rect 65258 4924 65566 4933
rect 65258 4922 65264 4924
rect 65320 4922 65344 4924
rect 65400 4922 65424 4924
rect 65480 4922 65504 4924
rect 65560 4922 65566 4924
rect 65320 4870 65322 4922
rect 65502 4870 65504 4922
rect 65258 4868 65264 4870
rect 65320 4868 65344 4870
rect 65400 4868 65424 4870
rect 65480 4868 65504 4870
rect 65560 4868 65566 4870
rect 65258 4859 65566 4868
rect 65628 4758 65656 5102
rect 65720 5030 65748 5782
rect 65708 5024 65760 5030
rect 65708 4966 65760 4972
rect 65616 4752 65668 4758
rect 65616 4694 65668 4700
rect 65156 4004 65208 4010
rect 65156 3946 65208 3952
rect 65258 3836 65566 3845
rect 65258 3834 65264 3836
rect 65320 3834 65344 3836
rect 65400 3834 65424 3836
rect 65480 3834 65504 3836
rect 65560 3834 65566 3836
rect 65320 3782 65322 3834
rect 65502 3782 65504 3834
rect 65258 3780 65264 3782
rect 65320 3780 65344 3782
rect 65400 3780 65424 3782
rect 65480 3780 65504 3782
rect 65560 3780 65566 3782
rect 65258 3771 65566 3780
rect 65156 3664 65208 3670
rect 65156 3606 65208 3612
rect 65064 2100 65116 2106
rect 65064 2042 65116 2048
rect 65168 1562 65196 3606
rect 65628 2922 65656 4694
rect 65616 2916 65668 2922
rect 65616 2858 65668 2864
rect 65258 2748 65566 2757
rect 65258 2746 65264 2748
rect 65320 2746 65344 2748
rect 65400 2746 65424 2748
rect 65480 2746 65504 2748
rect 65560 2746 65566 2748
rect 65320 2694 65322 2746
rect 65502 2694 65504 2746
rect 65258 2692 65264 2694
rect 65320 2692 65344 2694
rect 65400 2692 65424 2694
rect 65480 2692 65504 2694
rect 65560 2692 65566 2694
rect 65258 2683 65566 2692
rect 65720 2650 65748 4966
rect 65996 4826 66024 6190
rect 66088 5166 66116 7958
rect 66076 5160 66128 5166
rect 66076 5102 66128 5108
rect 65984 4820 66036 4826
rect 65984 4762 66036 4768
rect 65984 3936 66036 3942
rect 65984 3878 66036 3884
rect 65996 3466 66024 3878
rect 65984 3460 66036 3466
rect 65984 3402 66036 3408
rect 65800 3052 65852 3058
rect 65800 2994 65852 3000
rect 65708 2644 65760 2650
rect 65708 2586 65760 2592
rect 65248 2440 65300 2446
rect 65248 2382 65300 2388
rect 65260 1970 65288 2382
rect 65720 1970 65748 2586
rect 65248 1964 65300 1970
rect 65248 1906 65300 1912
rect 65708 1964 65760 1970
rect 65708 1906 65760 1912
rect 65812 1902 65840 2994
rect 65800 1896 65852 1902
rect 65800 1838 65852 1844
rect 65258 1660 65566 1669
rect 65258 1658 65264 1660
rect 65320 1658 65344 1660
rect 65400 1658 65424 1660
rect 65480 1658 65504 1660
rect 65560 1658 65566 1660
rect 65320 1606 65322 1658
rect 65502 1606 65504 1658
rect 65258 1604 65264 1606
rect 65320 1604 65344 1606
rect 65400 1604 65424 1606
rect 65480 1604 65504 1606
rect 65560 1604 65566 1606
rect 65258 1595 65566 1604
rect 65156 1556 65208 1562
rect 65156 1498 65208 1504
rect 64972 1012 65024 1018
rect 64972 954 65024 960
rect 65812 882 65840 1838
rect 65996 1358 66024 3402
rect 66180 2038 66208 11154
rect 66364 2582 66392 11222
rect 66456 3534 66484 16050
rect 66444 3528 66496 3534
rect 66444 3470 66496 3476
rect 66352 2576 66404 2582
rect 66352 2518 66404 2524
rect 66168 2032 66220 2038
rect 66168 1974 66220 1980
rect 65984 1352 66036 1358
rect 65984 1294 66036 1300
rect 65800 876 65852 882
rect 65800 818 65852 824
rect 65258 572 65566 581
rect 65258 570 65264 572
rect 65320 570 65344 572
rect 65400 570 65424 572
rect 65480 570 65504 572
rect 65560 570 65566 572
rect 65320 518 65322 570
rect 65502 518 65504 570
rect 65258 516 65264 518
rect 65320 516 65344 518
rect 65400 516 65424 518
rect 65480 516 65504 518
rect 65560 516 65566 518
rect 65258 507 65566 516
<< via2 >>
rect 35346 45056 35402 45112
rect 24858 44920 24914 44976
rect 12530 44648 12586 44704
rect 16210 44648 16266 44704
rect 2004 44634 2060 44636
rect 2084 44634 2140 44636
rect 2164 44634 2220 44636
rect 2244 44634 2300 44636
rect 2004 44582 2050 44634
rect 2050 44582 2060 44634
rect 2084 44582 2114 44634
rect 2114 44582 2126 44634
rect 2126 44582 2140 44634
rect 2164 44582 2178 44634
rect 2178 44582 2190 44634
rect 2190 44582 2220 44634
rect 2244 44582 2254 44634
rect 2254 44582 2300 44634
rect 2004 44580 2060 44582
rect 2084 44580 2140 44582
rect 2164 44580 2220 44582
rect 2244 44580 2300 44582
rect 6182 44532 6238 44568
rect 6182 44512 6184 44532
rect 6184 44512 6236 44532
rect 6236 44512 6238 44532
rect 6734 44532 6790 44568
rect 6734 44512 6736 44532
rect 6736 44512 6788 44532
rect 6788 44512 6790 44532
rect 7286 44532 7342 44568
rect 7286 44512 7288 44532
rect 7288 44512 7340 44532
rect 7340 44512 7342 44532
rect 7838 44532 7894 44568
rect 7838 44512 7840 44532
rect 7840 44512 7892 44532
rect 7892 44512 7894 44532
rect 8390 44532 8446 44568
rect 8390 44512 8392 44532
rect 8392 44512 8444 44532
rect 8444 44512 8446 44532
rect 8942 44532 8998 44568
rect 8942 44512 8944 44532
rect 8944 44512 8996 44532
rect 8996 44512 8998 44532
rect 9494 44532 9550 44568
rect 9494 44512 9496 44532
rect 9496 44512 9548 44532
rect 9548 44512 9550 44532
rect 10046 44532 10102 44568
rect 10046 44512 10048 44532
rect 10048 44512 10100 44532
rect 10100 44512 10102 44532
rect 10598 44532 10654 44568
rect 10598 44512 10600 44532
rect 10600 44512 10652 44532
rect 10652 44512 10654 44532
rect 12254 44532 12310 44568
rect 12254 44512 12256 44532
rect 12256 44512 12308 44532
rect 12308 44512 12310 44532
rect 12806 44532 12862 44568
rect 12806 44512 12808 44532
rect 12808 44512 12860 44532
rect 12860 44512 12862 44532
rect 13542 44532 13598 44568
rect 13542 44512 13544 44532
rect 13544 44512 13596 44532
rect 13596 44512 13598 44532
rect 13818 44532 13874 44568
rect 13818 44512 13820 44532
rect 13820 44512 13872 44532
rect 13872 44512 13874 44532
rect 15474 44532 15530 44568
rect 15474 44512 15476 44532
rect 15476 44512 15528 44532
rect 15528 44512 15530 44532
rect 15934 44532 15990 44568
rect 15934 44512 15936 44532
rect 15936 44512 15988 44532
rect 15988 44512 15990 44532
rect 16670 44532 16726 44568
rect 16670 44512 16672 44532
rect 16672 44512 16724 44532
rect 16724 44512 16726 44532
rect 17222 44648 17278 44704
rect 16946 44532 17002 44568
rect 16946 44512 16948 44532
rect 16948 44512 17000 44532
rect 17000 44512 17002 44532
rect 2924 44090 2980 44092
rect 3004 44090 3060 44092
rect 3084 44090 3140 44092
rect 3164 44090 3220 44092
rect 2924 44038 2970 44090
rect 2970 44038 2980 44090
rect 3004 44038 3034 44090
rect 3034 44038 3046 44090
rect 3046 44038 3060 44090
rect 3084 44038 3098 44090
rect 3098 44038 3110 44090
rect 3110 44038 3140 44090
rect 3164 44038 3174 44090
rect 3174 44038 3220 44090
rect 2924 44036 2980 44038
rect 3004 44036 3060 44038
rect 3084 44036 3140 44038
rect 3164 44036 3220 44038
rect 2004 43546 2060 43548
rect 2084 43546 2140 43548
rect 2164 43546 2220 43548
rect 2244 43546 2300 43548
rect 2004 43494 2050 43546
rect 2050 43494 2060 43546
rect 2084 43494 2114 43546
rect 2114 43494 2126 43546
rect 2126 43494 2140 43546
rect 2164 43494 2178 43546
rect 2178 43494 2190 43546
rect 2190 43494 2220 43546
rect 2244 43494 2254 43546
rect 2254 43494 2300 43546
rect 2004 43492 2060 43494
rect 2084 43492 2140 43494
rect 2164 43492 2220 43494
rect 2244 43492 2300 43494
rect 11150 43852 11206 43888
rect 11150 43832 11152 43852
rect 11152 43832 11204 43852
rect 11204 43832 11206 43852
rect 2924 43002 2980 43004
rect 3004 43002 3060 43004
rect 3084 43002 3140 43004
rect 3164 43002 3220 43004
rect 2924 42950 2970 43002
rect 2970 42950 2980 43002
rect 3004 42950 3034 43002
rect 3034 42950 3046 43002
rect 3046 42950 3060 43002
rect 3084 42950 3098 43002
rect 3098 42950 3110 43002
rect 3110 42950 3140 43002
rect 3164 42950 3174 43002
rect 3174 42950 3220 43002
rect 2924 42948 2980 42950
rect 3004 42948 3060 42950
rect 3084 42948 3140 42950
rect 3164 42948 3220 42950
rect 2004 42458 2060 42460
rect 2084 42458 2140 42460
rect 2164 42458 2220 42460
rect 2244 42458 2300 42460
rect 2004 42406 2050 42458
rect 2050 42406 2060 42458
rect 2084 42406 2114 42458
rect 2114 42406 2126 42458
rect 2126 42406 2140 42458
rect 2164 42406 2178 42458
rect 2178 42406 2190 42458
rect 2190 42406 2220 42458
rect 2244 42406 2254 42458
rect 2254 42406 2300 42458
rect 2004 42404 2060 42406
rect 2084 42404 2140 42406
rect 2164 42404 2220 42406
rect 2244 42404 2300 42406
rect 2924 41914 2980 41916
rect 3004 41914 3060 41916
rect 3084 41914 3140 41916
rect 3164 41914 3220 41916
rect 2924 41862 2970 41914
rect 2970 41862 2980 41914
rect 3004 41862 3034 41914
rect 3034 41862 3046 41914
rect 3046 41862 3060 41914
rect 3084 41862 3098 41914
rect 3098 41862 3110 41914
rect 3110 41862 3140 41914
rect 3164 41862 3174 41914
rect 3174 41862 3220 41914
rect 2924 41860 2980 41862
rect 3004 41860 3060 41862
rect 3084 41860 3140 41862
rect 3164 41860 3220 41862
rect 2004 41370 2060 41372
rect 2084 41370 2140 41372
rect 2164 41370 2220 41372
rect 2244 41370 2300 41372
rect 2004 41318 2050 41370
rect 2050 41318 2060 41370
rect 2084 41318 2114 41370
rect 2114 41318 2126 41370
rect 2126 41318 2140 41370
rect 2164 41318 2178 41370
rect 2178 41318 2190 41370
rect 2190 41318 2220 41370
rect 2244 41318 2254 41370
rect 2254 41318 2300 41370
rect 2004 41316 2060 41318
rect 2084 41316 2140 41318
rect 2164 41316 2220 41318
rect 2244 41316 2300 41318
rect 2924 40826 2980 40828
rect 3004 40826 3060 40828
rect 3084 40826 3140 40828
rect 3164 40826 3220 40828
rect 2924 40774 2970 40826
rect 2970 40774 2980 40826
rect 3004 40774 3034 40826
rect 3034 40774 3046 40826
rect 3046 40774 3060 40826
rect 3084 40774 3098 40826
rect 3098 40774 3110 40826
rect 3110 40774 3140 40826
rect 3164 40774 3174 40826
rect 3174 40774 3220 40826
rect 2924 40772 2980 40774
rect 3004 40772 3060 40774
rect 3084 40772 3140 40774
rect 3164 40772 3220 40774
rect 2004 40282 2060 40284
rect 2084 40282 2140 40284
rect 2164 40282 2220 40284
rect 2244 40282 2300 40284
rect 2004 40230 2050 40282
rect 2050 40230 2060 40282
rect 2084 40230 2114 40282
rect 2114 40230 2126 40282
rect 2126 40230 2140 40282
rect 2164 40230 2178 40282
rect 2178 40230 2190 40282
rect 2190 40230 2220 40282
rect 2244 40230 2254 40282
rect 2254 40230 2300 40282
rect 2004 40228 2060 40230
rect 2084 40228 2140 40230
rect 2164 40228 2220 40230
rect 2244 40228 2300 40230
rect 2924 39738 2980 39740
rect 3004 39738 3060 39740
rect 3084 39738 3140 39740
rect 3164 39738 3220 39740
rect 2924 39686 2970 39738
rect 2970 39686 2980 39738
rect 3004 39686 3034 39738
rect 3034 39686 3046 39738
rect 3046 39686 3060 39738
rect 3084 39686 3098 39738
rect 3098 39686 3110 39738
rect 3110 39686 3140 39738
rect 3164 39686 3174 39738
rect 3174 39686 3220 39738
rect 2924 39684 2980 39686
rect 3004 39684 3060 39686
rect 3084 39684 3140 39686
rect 3164 39684 3220 39686
rect 2004 39194 2060 39196
rect 2084 39194 2140 39196
rect 2164 39194 2220 39196
rect 2244 39194 2300 39196
rect 2004 39142 2050 39194
rect 2050 39142 2060 39194
rect 2084 39142 2114 39194
rect 2114 39142 2126 39194
rect 2126 39142 2140 39194
rect 2164 39142 2178 39194
rect 2178 39142 2190 39194
rect 2190 39142 2220 39194
rect 2244 39142 2254 39194
rect 2254 39142 2300 39194
rect 2004 39140 2060 39142
rect 2084 39140 2140 39142
rect 2164 39140 2220 39142
rect 2244 39140 2300 39142
rect 2924 38650 2980 38652
rect 3004 38650 3060 38652
rect 3084 38650 3140 38652
rect 3164 38650 3220 38652
rect 2924 38598 2970 38650
rect 2970 38598 2980 38650
rect 3004 38598 3034 38650
rect 3034 38598 3046 38650
rect 3046 38598 3060 38650
rect 3084 38598 3098 38650
rect 3098 38598 3110 38650
rect 3110 38598 3140 38650
rect 3164 38598 3174 38650
rect 3174 38598 3220 38650
rect 2924 38596 2980 38598
rect 3004 38596 3060 38598
rect 3084 38596 3140 38598
rect 3164 38596 3220 38598
rect 2004 38106 2060 38108
rect 2084 38106 2140 38108
rect 2164 38106 2220 38108
rect 2244 38106 2300 38108
rect 2004 38054 2050 38106
rect 2050 38054 2060 38106
rect 2084 38054 2114 38106
rect 2114 38054 2126 38106
rect 2126 38054 2140 38106
rect 2164 38054 2178 38106
rect 2178 38054 2190 38106
rect 2190 38054 2220 38106
rect 2244 38054 2254 38106
rect 2254 38054 2300 38106
rect 2004 38052 2060 38054
rect 2084 38052 2140 38054
rect 2164 38052 2220 38054
rect 2244 38052 2300 38054
rect 2924 37562 2980 37564
rect 3004 37562 3060 37564
rect 3084 37562 3140 37564
rect 3164 37562 3220 37564
rect 2924 37510 2970 37562
rect 2970 37510 2980 37562
rect 3004 37510 3034 37562
rect 3034 37510 3046 37562
rect 3046 37510 3060 37562
rect 3084 37510 3098 37562
rect 3098 37510 3110 37562
rect 3110 37510 3140 37562
rect 3164 37510 3174 37562
rect 3174 37510 3220 37562
rect 2924 37508 2980 37510
rect 3004 37508 3060 37510
rect 3084 37508 3140 37510
rect 3164 37508 3220 37510
rect 11426 40588 11482 40624
rect 11426 40568 11428 40588
rect 11428 40568 11480 40588
rect 11480 40568 11482 40588
rect 11610 39616 11666 39672
rect 15290 43852 15346 43888
rect 15290 43832 15292 43852
rect 15292 43832 15344 43852
rect 15344 43832 15346 43852
rect 12714 39888 12770 39944
rect 12070 38412 12126 38448
rect 12070 38392 12072 38412
rect 12072 38392 12124 38412
rect 12124 38392 12126 38412
rect 2004 37018 2060 37020
rect 2084 37018 2140 37020
rect 2164 37018 2220 37020
rect 2244 37018 2300 37020
rect 2004 36966 2050 37018
rect 2050 36966 2060 37018
rect 2084 36966 2114 37018
rect 2114 36966 2126 37018
rect 2126 36966 2140 37018
rect 2164 36966 2178 37018
rect 2178 36966 2190 37018
rect 2190 36966 2220 37018
rect 2244 36966 2254 37018
rect 2254 36966 2300 37018
rect 2004 36964 2060 36966
rect 2084 36964 2140 36966
rect 2164 36964 2220 36966
rect 2244 36964 2300 36966
rect 15658 41268 15714 41304
rect 15658 41248 15660 41268
rect 15660 41248 15712 41268
rect 15712 41248 15714 41268
rect 16854 42200 16910 42256
rect 17958 43716 18014 43752
rect 17958 43696 17960 43716
rect 17960 43696 18012 43716
rect 18012 43696 18014 43716
rect 18786 43424 18842 43480
rect 19798 43732 19800 43752
rect 19800 43732 19852 43752
rect 19852 43732 19854 43752
rect 19798 43696 19854 43732
rect 14830 37712 14886 37768
rect 12162 35944 12218 36000
rect 8206 35708 8208 35728
rect 8208 35708 8260 35728
rect 8260 35708 8262 35728
rect 8206 35672 8262 35708
rect 15106 37304 15162 37360
rect 15106 36624 15162 36680
rect 19154 41384 19210 41440
rect 19522 38664 19578 38720
rect 19522 37032 19578 37088
rect 15290 36624 15346 36680
rect 20902 40840 20958 40896
rect 26606 44648 26662 44704
rect 26238 44376 26294 44432
rect 22374 41520 22430 41576
rect 24030 41656 24086 41712
rect 21638 37168 21694 37224
rect 20350 36896 20406 36952
rect 21638 36896 21694 36952
rect 23202 36760 23258 36816
rect 19706 35944 19762 36000
rect 26790 44396 26846 44432
rect 26790 44376 26792 44396
rect 26792 44376 26844 44396
rect 26844 44376 26846 44396
rect 27526 44396 27582 44432
rect 27526 44376 27528 44396
rect 27528 44376 27580 44396
rect 27580 44376 27582 44396
rect 26514 43696 26570 43752
rect 26606 42628 26662 42664
rect 26606 42608 26608 42628
rect 26608 42608 26660 42628
rect 26660 42608 26662 42628
rect 24858 40568 24914 40624
rect 25502 40976 25558 41032
rect 24122 38664 24178 38720
rect 25134 38548 25190 38584
rect 25134 38528 25136 38548
rect 25136 38528 25188 38548
rect 25188 38528 25190 38548
rect 22006 35808 22062 35864
rect 24030 36216 24086 36272
rect 24766 36760 24822 36816
rect 26146 41248 26202 41304
rect 25962 40704 26018 40760
rect 27066 41928 27122 41984
rect 25962 39344 26018 39400
rect 25686 38700 25688 38720
rect 25688 38700 25740 38720
rect 25740 38700 25742 38720
rect 25686 38664 25742 38700
rect 26146 38528 26202 38584
rect 27802 42628 27858 42664
rect 27802 42608 27804 42628
rect 27804 42608 27856 42628
rect 27856 42608 27858 42628
rect 27710 41928 27766 41984
rect 27158 41112 27214 41168
rect 27066 40568 27122 40624
rect 26054 37032 26110 37088
rect 25502 36080 25558 36136
rect 23570 35808 23626 35864
rect 24490 35808 24546 35864
rect 24766 35844 24768 35864
rect 24768 35844 24820 35864
rect 24820 35844 24822 35864
rect 24766 35808 24822 35844
rect 27710 41384 27766 41440
rect 31758 44784 31814 44840
rect 28722 41792 28778 41848
rect 27710 40296 27766 40352
rect 27802 38820 27858 38856
rect 27802 38800 27804 38820
rect 27804 38800 27856 38820
rect 27856 38800 27858 38820
rect 27618 38392 27674 38448
rect 27894 37304 27950 37360
rect 28538 37304 28594 37360
rect 25870 35808 25926 35864
rect 29642 43308 29698 43344
rect 29642 43288 29644 43308
rect 29644 43288 29696 43308
rect 29696 43288 29698 43308
rect 29274 40468 29276 40488
rect 29276 40468 29328 40488
rect 29328 40468 29330 40488
rect 29274 40432 29330 40468
rect 28814 39616 28870 39672
rect 29090 39480 29146 39536
rect 29734 40160 29790 40216
rect 29642 39480 29698 39536
rect 29458 38800 29514 38856
rect 29550 38276 29606 38312
rect 29550 38256 29552 38276
rect 29552 38256 29604 38276
rect 29604 38256 29606 38276
rect 29090 37032 29146 37088
rect 28998 36216 29054 36272
rect 15014 35672 15070 35728
rect 20074 35672 20130 35728
rect 21362 35672 21418 35728
rect 22190 35692 22246 35728
rect 22190 35672 22192 35692
rect 22192 35672 22244 35692
rect 22244 35672 22246 35692
rect 23018 35672 23074 35728
rect 23202 35672 23258 35728
rect 25226 35672 25282 35728
rect 30102 36488 30158 36544
rect 30010 35808 30066 35864
rect 30562 43424 30618 43480
rect 30378 41964 30380 41984
rect 30380 41964 30432 41984
rect 30432 41964 30434 41984
rect 30378 41928 30434 41964
rect 30378 40976 30434 41032
rect 31390 43732 31392 43752
rect 31392 43732 31444 43752
rect 31444 43732 31446 43752
rect 31390 43696 31446 43732
rect 31206 43288 31262 43344
rect 31666 43424 31722 43480
rect 31114 41928 31170 41984
rect 31114 41656 31170 41712
rect 30838 39480 30894 39536
rect 31206 40468 31208 40488
rect 31208 40468 31260 40488
rect 31260 40468 31262 40488
rect 31206 40432 31262 40468
rect 31666 40588 31722 40624
rect 31666 40568 31668 40588
rect 31668 40568 31720 40588
rect 31720 40568 31722 40588
rect 31206 38700 31208 38720
rect 31208 38700 31260 38720
rect 31260 38700 31262 38720
rect 31206 38664 31262 38700
rect 30378 36760 30434 36816
rect 30194 35808 30250 35864
rect 30470 36352 30526 36408
rect 31850 42608 31906 42664
rect 31850 41540 31906 41576
rect 31850 41520 31852 41540
rect 31852 41520 31904 41540
rect 31904 41520 31906 41540
rect 31850 40996 31906 41032
rect 31850 40976 31852 40996
rect 31852 40976 31904 40996
rect 31904 40976 31906 40996
rect 32494 42472 32550 42528
rect 32034 40024 32090 40080
rect 33046 42200 33102 42256
rect 33506 42200 33562 42256
rect 32862 39752 32918 39808
rect 32494 39208 32550 39264
rect 32494 38800 32550 38856
rect 32678 39244 32680 39264
rect 32680 39244 32732 39264
rect 32732 39244 32734 39264
rect 32678 39208 32734 39244
rect 32770 39072 32826 39128
rect 32402 37168 32458 37224
rect 32954 39344 33010 39400
rect 33138 37848 33194 37904
rect 32862 36352 32918 36408
rect 31666 35944 31722 36000
rect 34518 41420 34520 41440
rect 34520 41420 34572 41440
rect 34572 41420 34574 41440
rect 34518 41384 34574 41420
rect 35070 42356 35126 42392
rect 35070 42336 35072 42356
rect 35072 42336 35124 42356
rect 35124 42336 35126 42356
rect 34794 41112 34850 41168
rect 34150 38256 34206 38312
rect 33690 37304 33746 37360
rect 33414 35944 33470 36000
rect 31114 35808 31170 35864
rect 33046 35808 33102 35864
rect 34426 38256 34482 38312
rect 34334 38120 34390 38176
rect 34518 37460 34574 37496
rect 34518 37440 34520 37460
rect 34520 37440 34572 37460
rect 34572 37440 34574 37460
rect 34426 37168 34482 37224
rect 35254 39480 35310 39536
rect 36818 43016 36874 43072
rect 35806 40160 35862 40216
rect 36450 40840 36506 40896
rect 36634 41520 36690 41576
rect 51004 44634 51060 44636
rect 51084 44634 51140 44636
rect 51164 44634 51220 44636
rect 51244 44634 51300 44636
rect 51004 44582 51050 44634
rect 51050 44582 51060 44634
rect 51084 44582 51114 44634
rect 51114 44582 51126 44634
rect 51126 44582 51140 44634
rect 51164 44582 51178 44634
rect 51178 44582 51190 44634
rect 51190 44582 51220 44634
rect 51244 44582 51254 44634
rect 51254 44582 51300 44634
rect 51004 44580 51060 44582
rect 51084 44580 51140 44582
rect 51164 44580 51220 44582
rect 51244 44580 51300 44582
rect 37094 41268 37150 41304
rect 37094 41248 37096 41268
rect 37096 41248 37148 41268
rect 37148 41248 37150 41268
rect 37002 41112 37058 41168
rect 37094 40996 37150 41032
rect 37094 40976 37096 40996
rect 37096 40976 37148 40996
rect 37148 40976 37150 40996
rect 35806 37304 35862 37360
rect 37278 40296 37334 40352
rect 37370 40024 37426 40080
rect 36818 36896 36874 36952
rect 38014 37984 38070 38040
rect 38658 39752 38714 39808
rect 38658 39208 38714 39264
rect 38934 37984 38990 38040
rect 41878 41928 41934 41984
rect 40774 38800 40830 38856
rect 41694 38820 41750 38856
rect 41694 38800 41696 38820
rect 41696 38800 41748 38820
rect 41748 38800 41750 38820
rect 44822 41792 44878 41848
rect 45558 42064 45614 42120
rect 43626 38800 43682 38856
rect 44546 38800 44602 38856
rect 45190 39616 45246 39672
rect 45466 39616 45522 39672
rect 46662 38820 46718 38856
rect 46662 38800 46664 38820
rect 46664 38800 46716 38820
rect 46716 38800 46718 38820
rect 47490 38820 47546 38856
rect 47490 38800 47492 38820
rect 47492 38800 47544 38820
rect 47544 38800 47546 38820
rect 43810 37612 43812 37632
rect 43812 37612 43864 37632
rect 43864 37612 43866 37632
rect 43810 37576 43866 37612
rect 51924 44090 51980 44092
rect 52004 44090 52060 44092
rect 52084 44090 52140 44092
rect 52164 44090 52220 44092
rect 51924 44038 51970 44090
rect 51970 44038 51980 44090
rect 52004 44038 52034 44090
rect 52034 44038 52046 44090
rect 52046 44038 52060 44090
rect 52084 44038 52098 44090
rect 52098 44038 52110 44090
rect 52110 44038 52140 44090
rect 52164 44038 52174 44090
rect 52174 44038 52220 44090
rect 51924 44036 51980 44038
rect 52004 44036 52060 44038
rect 52084 44036 52140 44038
rect 52164 44036 52220 44038
rect 51004 43546 51060 43548
rect 51084 43546 51140 43548
rect 51164 43546 51220 43548
rect 51244 43546 51300 43548
rect 51004 43494 51050 43546
rect 51050 43494 51060 43546
rect 51084 43494 51114 43546
rect 51114 43494 51126 43546
rect 51126 43494 51140 43546
rect 51164 43494 51178 43546
rect 51178 43494 51190 43546
rect 51190 43494 51220 43546
rect 51244 43494 51254 43546
rect 51254 43494 51300 43546
rect 51004 43492 51060 43494
rect 51084 43492 51140 43494
rect 51164 43492 51220 43494
rect 51244 43492 51300 43494
rect 51004 42458 51060 42460
rect 51084 42458 51140 42460
rect 51164 42458 51220 42460
rect 51244 42458 51300 42460
rect 51004 42406 51050 42458
rect 51050 42406 51060 42458
rect 51084 42406 51114 42458
rect 51114 42406 51126 42458
rect 51126 42406 51140 42458
rect 51164 42406 51178 42458
rect 51178 42406 51190 42458
rect 51190 42406 51220 42458
rect 51244 42406 51254 42458
rect 51254 42406 51300 42458
rect 51004 42404 51060 42406
rect 51084 42404 51140 42406
rect 51164 42404 51220 42406
rect 51244 42404 51300 42406
rect 51924 43002 51980 43004
rect 52004 43002 52060 43004
rect 52084 43002 52140 43004
rect 52164 43002 52220 43004
rect 51924 42950 51970 43002
rect 51970 42950 51980 43002
rect 52004 42950 52034 43002
rect 52034 42950 52046 43002
rect 52046 42950 52060 43002
rect 52084 42950 52098 43002
rect 52098 42950 52110 43002
rect 52110 42950 52140 43002
rect 52164 42950 52174 43002
rect 52174 42950 52220 43002
rect 51924 42948 51980 42950
rect 52004 42948 52060 42950
rect 52084 42948 52140 42950
rect 52164 42948 52220 42950
rect 51924 41914 51980 41916
rect 52004 41914 52060 41916
rect 52084 41914 52140 41916
rect 52164 41914 52220 41916
rect 51924 41862 51970 41914
rect 51970 41862 51980 41914
rect 52004 41862 52034 41914
rect 52034 41862 52046 41914
rect 52046 41862 52060 41914
rect 52084 41862 52098 41914
rect 52098 41862 52110 41914
rect 52110 41862 52140 41914
rect 52164 41862 52174 41914
rect 52174 41862 52220 41914
rect 51924 41860 51980 41862
rect 52004 41860 52060 41862
rect 52084 41860 52140 41862
rect 52164 41860 52220 41862
rect 49054 40704 49110 40760
rect 49146 39616 49202 39672
rect 50618 40840 50674 40896
rect 50526 39636 50582 39672
rect 50526 39616 50528 39636
rect 50528 39616 50580 39636
rect 50580 39616 50582 39636
rect 50066 37848 50122 37904
rect 51004 41370 51060 41372
rect 51084 41370 51140 41372
rect 51164 41370 51220 41372
rect 51244 41370 51300 41372
rect 51004 41318 51050 41370
rect 51050 41318 51060 41370
rect 51084 41318 51114 41370
rect 51114 41318 51126 41370
rect 51126 41318 51140 41370
rect 51164 41318 51178 41370
rect 51178 41318 51190 41370
rect 51190 41318 51220 41370
rect 51244 41318 51254 41370
rect 51254 41318 51300 41370
rect 51004 41316 51060 41318
rect 51084 41316 51140 41318
rect 51164 41316 51220 41318
rect 51244 41316 51300 41318
rect 51924 40826 51980 40828
rect 52004 40826 52060 40828
rect 52084 40826 52140 40828
rect 52164 40826 52220 40828
rect 51924 40774 51970 40826
rect 51970 40774 51980 40826
rect 52004 40774 52034 40826
rect 52034 40774 52046 40826
rect 52046 40774 52060 40826
rect 52084 40774 52098 40826
rect 52098 40774 52110 40826
rect 52110 40774 52140 40826
rect 52164 40774 52174 40826
rect 52174 40774 52220 40826
rect 51924 40772 51980 40774
rect 52004 40772 52060 40774
rect 52084 40772 52140 40774
rect 52164 40772 52220 40774
rect 51004 40282 51060 40284
rect 51084 40282 51140 40284
rect 51164 40282 51220 40284
rect 51244 40282 51300 40284
rect 51004 40230 51050 40282
rect 51050 40230 51060 40282
rect 51084 40230 51114 40282
rect 51114 40230 51126 40282
rect 51126 40230 51140 40282
rect 51164 40230 51178 40282
rect 51178 40230 51190 40282
rect 51190 40230 51220 40282
rect 51244 40230 51254 40282
rect 51254 40230 51300 40282
rect 51004 40228 51060 40230
rect 51084 40228 51140 40230
rect 51164 40228 51220 40230
rect 51244 40228 51300 40230
rect 51924 39738 51980 39740
rect 52004 39738 52060 39740
rect 52084 39738 52140 39740
rect 52164 39738 52220 39740
rect 51924 39686 51970 39738
rect 51970 39686 51980 39738
rect 52004 39686 52034 39738
rect 52034 39686 52046 39738
rect 52046 39686 52060 39738
rect 52084 39686 52098 39738
rect 52098 39686 52110 39738
rect 52110 39686 52140 39738
rect 52164 39686 52174 39738
rect 52174 39686 52220 39738
rect 51924 39684 51980 39686
rect 52004 39684 52060 39686
rect 52084 39684 52140 39686
rect 52164 39684 52220 39686
rect 51004 39194 51060 39196
rect 51084 39194 51140 39196
rect 51164 39194 51220 39196
rect 51244 39194 51300 39196
rect 51004 39142 51050 39194
rect 51050 39142 51060 39194
rect 51084 39142 51114 39194
rect 51114 39142 51126 39194
rect 51126 39142 51140 39194
rect 51164 39142 51178 39194
rect 51178 39142 51190 39194
rect 51190 39142 51220 39194
rect 51244 39142 51254 39194
rect 51254 39142 51300 39194
rect 51004 39140 51060 39142
rect 51084 39140 51140 39142
rect 51164 39140 51220 39142
rect 51244 39140 51300 39142
rect 51924 38650 51980 38652
rect 52004 38650 52060 38652
rect 52084 38650 52140 38652
rect 52164 38650 52220 38652
rect 51924 38598 51970 38650
rect 51970 38598 51980 38650
rect 52004 38598 52034 38650
rect 52034 38598 52046 38650
rect 52046 38598 52060 38650
rect 52084 38598 52098 38650
rect 52098 38598 52110 38650
rect 52110 38598 52140 38650
rect 52164 38598 52174 38650
rect 52174 38598 52220 38650
rect 51924 38596 51980 38598
rect 52004 38596 52060 38598
rect 52084 38596 52140 38598
rect 52164 38596 52220 38598
rect 51004 38106 51060 38108
rect 51084 38106 51140 38108
rect 51164 38106 51220 38108
rect 51244 38106 51300 38108
rect 51004 38054 51050 38106
rect 51050 38054 51060 38106
rect 51084 38054 51114 38106
rect 51114 38054 51126 38106
rect 51126 38054 51140 38106
rect 51164 38054 51178 38106
rect 51178 38054 51190 38106
rect 51190 38054 51220 38106
rect 51244 38054 51254 38106
rect 51254 38054 51300 38106
rect 51004 38052 51060 38054
rect 51084 38052 51140 38054
rect 51164 38052 51220 38054
rect 51244 38052 51300 38054
rect 51924 37562 51980 37564
rect 52004 37562 52060 37564
rect 52084 37562 52140 37564
rect 52164 37562 52220 37564
rect 51924 37510 51970 37562
rect 51970 37510 51980 37562
rect 52004 37510 52034 37562
rect 52034 37510 52046 37562
rect 52046 37510 52060 37562
rect 52084 37510 52098 37562
rect 52098 37510 52110 37562
rect 52110 37510 52140 37562
rect 52164 37510 52174 37562
rect 52174 37510 52220 37562
rect 51924 37508 51980 37510
rect 52004 37508 52060 37510
rect 52084 37508 52140 37510
rect 52164 37508 52220 37510
rect 52826 38936 52882 38992
rect 51004 37018 51060 37020
rect 51084 37018 51140 37020
rect 51164 37018 51220 37020
rect 51244 37018 51300 37020
rect 51004 36966 51050 37018
rect 51050 36966 51060 37018
rect 51084 36966 51114 37018
rect 51114 36966 51126 37018
rect 51126 36966 51140 37018
rect 51164 36966 51178 37018
rect 51178 36966 51190 37018
rect 51190 36966 51220 37018
rect 51244 36966 51254 37018
rect 51254 36966 51300 37018
rect 51004 36964 51060 36966
rect 51084 36964 51140 36966
rect 51164 36964 51220 36966
rect 51244 36964 51300 36966
rect 57058 40568 57114 40624
rect 55402 37732 55458 37768
rect 55402 37712 55404 37732
rect 55404 37712 55456 37732
rect 55456 37712 55458 37732
rect 55862 37732 55918 37768
rect 55862 37712 55864 37732
rect 55864 37712 55916 37732
rect 55916 37712 55918 37732
rect 57702 39924 57704 39944
rect 57704 39924 57756 39944
rect 57756 39924 57758 39944
rect 57702 39888 57758 39924
rect 60738 42608 60794 42664
rect 62854 40976 62910 41032
rect 60738 40160 60794 40216
rect 62026 37304 62082 37360
rect 37278 36216 37334 36272
rect 34426 36080 34482 36136
rect 34518 35808 34574 35864
rect 38566 35808 38622 35864
rect 30286 35672 30342 35728
rect 30470 35672 30526 35728
rect 36542 35672 36598 35728
rect 38658 35672 38714 35728
rect 42706 35808 42762 35864
rect 56414 35672 56470 35728
rect 62118 35944 62174 36000
rect 62578 36216 62634 36272
rect 62670 36080 62726 36136
rect 62670 31184 62726 31240
rect 48962 1808 49018 1864
rect 49238 1808 49294 1864
rect 49698 1844 49700 1864
rect 49700 1844 49752 1864
rect 49752 1844 49754 1864
rect 49698 1808 49754 1844
rect 63222 38256 63278 38312
rect 63590 36252 63592 36272
rect 63592 36252 63644 36272
rect 63644 36252 63646 36272
rect 63590 36216 63646 36252
rect 63498 34720 63554 34776
rect 63682 34584 63738 34640
rect 64344 37018 64400 37020
rect 64424 37018 64480 37020
rect 64504 37018 64560 37020
rect 64584 37018 64640 37020
rect 64344 36966 64390 37018
rect 64390 36966 64400 37018
rect 64424 36966 64454 37018
rect 64454 36966 64466 37018
rect 64466 36966 64480 37018
rect 64504 36966 64518 37018
rect 64518 36966 64530 37018
rect 64530 36966 64560 37018
rect 64584 36966 64594 37018
rect 64594 36966 64640 37018
rect 64344 36964 64400 36966
rect 64424 36964 64480 36966
rect 64504 36964 64560 36966
rect 64584 36964 64640 36966
rect 64344 35930 64400 35932
rect 64424 35930 64480 35932
rect 64504 35930 64560 35932
rect 64584 35930 64640 35932
rect 64344 35878 64390 35930
rect 64390 35878 64400 35930
rect 64424 35878 64454 35930
rect 64454 35878 64466 35930
rect 64466 35878 64480 35930
rect 64504 35878 64518 35930
rect 64518 35878 64530 35930
rect 64530 35878 64560 35930
rect 64584 35878 64594 35930
rect 64594 35878 64640 35930
rect 64344 35876 64400 35878
rect 64424 35876 64480 35878
rect 64504 35876 64560 35878
rect 64584 35876 64640 35878
rect 63958 35672 64014 35728
rect 64344 34842 64400 34844
rect 64424 34842 64480 34844
rect 64504 34842 64560 34844
rect 64584 34842 64640 34844
rect 64344 34790 64390 34842
rect 64390 34790 64400 34842
rect 64424 34790 64454 34842
rect 64454 34790 64466 34842
rect 64466 34790 64480 34842
rect 64504 34790 64518 34842
rect 64518 34790 64530 34842
rect 64530 34790 64560 34842
rect 64584 34790 64594 34842
rect 64594 34790 64640 34842
rect 64344 34788 64400 34790
rect 64424 34788 64480 34790
rect 64504 34788 64560 34790
rect 64584 34788 64640 34790
rect 64344 33754 64400 33756
rect 64424 33754 64480 33756
rect 64504 33754 64560 33756
rect 64584 33754 64640 33756
rect 64344 33702 64390 33754
rect 64390 33702 64400 33754
rect 64424 33702 64454 33754
rect 64454 33702 64466 33754
rect 64466 33702 64480 33754
rect 64504 33702 64518 33754
rect 64518 33702 64530 33754
rect 64530 33702 64560 33754
rect 64584 33702 64594 33754
rect 64594 33702 64640 33754
rect 64344 33700 64400 33702
rect 64424 33700 64480 33702
rect 64504 33700 64560 33702
rect 64584 33700 64640 33702
rect 64344 32666 64400 32668
rect 64424 32666 64480 32668
rect 64504 32666 64560 32668
rect 64584 32666 64640 32668
rect 64344 32614 64390 32666
rect 64390 32614 64400 32666
rect 64424 32614 64454 32666
rect 64454 32614 64466 32666
rect 64466 32614 64480 32666
rect 64504 32614 64518 32666
rect 64518 32614 64530 32666
rect 64530 32614 64560 32666
rect 64584 32614 64594 32666
rect 64594 32614 64640 32666
rect 64344 32612 64400 32614
rect 64424 32612 64480 32614
rect 64504 32612 64560 32614
rect 64584 32612 64640 32614
rect 65264 37562 65320 37564
rect 65344 37562 65400 37564
rect 65424 37562 65480 37564
rect 65504 37562 65560 37564
rect 65264 37510 65310 37562
rect 65310 37510 65320 37562
rect 65344 37510 65374 37562
rect 65374 37510 65386 37562
rect 65386 37510 65400 37562
rect 65424 37510 65438 37562
rect 65438 37510 65450 37562
rect 65450 37510 65480 37562
rect 65504 37510 65514 37562
rect 65514 37510 65560 37562
rect 65264 37508 65320 37510
rect 65344 37508 65400 37510
rect 65424 37508 65480 37510
rect 65504 37508 65560 37510
rect 65264 36474 65320 36476
rect 65344 36474 65400 36476
rect 65424 36474 65480 36476
rect 65504 36474 65560 36476
rect 65264 36422 65310 36474
rect 65310 36422 65320 36474
rect 65344 36422 65374 36474
rect 65374 36422 65386 36474
rect 65386 36422 65400 36474
rect 65424 36422 65438 36474
rect 65438 36422 65450 36474
rect 65450 36422 65480 36474
rect 65504 36422 65514 36474
rect 65514 36422 65560 36474
rect 65264 36420 65320 36422
rect 65344 36420 65400 36422
rect 65424 36420 65480 36422
rect 65504 36420 65560 36422
rect 65264 35386 65320 35388
rect 65344 35386 65400 35388
rect 65424 35386 65480 35388
rect 65504 35386 65560 35388
rect 65264 35334 65310 35386
rect 65310 35334 65320 35386
rect 65344 35334 65374 35386
rect 65374 35334 65386 35386
rect 65386 35334 65400 35386
rect 65424 35334 65438 35386
rect 65438 35334 65450 35386
rect 65450 35334 65480 35386
rect 65504 35334 65514 35386
rect 65514 35334 65560 35386
rect 65264 35332 65320 35334
rect 65344 35332 65400 35334
rect 65424 35332 65480 35334
rect 65504 35332 65560 35334
rect 65264 34298 65320 34300
rect 65344 34298 65400 34300
rect 65424 34298 65480 34300
rect 65504 34298 65560 34300
rect 65264 34246 65310 34298
rect 65310 34246 65320 34298
rect 65344 34246 65374 34298
rect 65374 34246 65386 34298
rect 65386 34246 65400 34298
rect 65424 34246 65438 34298
rect 65438 34246 65450 34298
rect 65450 34246 65480 34298
rect 65504 34246 65514 34298
rect 65514 34246 65560 34298
rect 65264 34244 65320 34246
rect 65344 34244 65400 34246
rect 65424 34244 65480 34246
rect 65504 34244 65560 34246
rect 64344 31578 64400 31580
rect 64424 31578 64480 31580
rect 64504 31578 64560 31580
rect 64584 31578 64640 31580
rect 64344 31526 64390 31578
rect 64390 31526 64400 31578
rect 64424 31526 64454 31578
rect 64454 31526 64466 31578
rect 64466 31526 64480 31578
rect 64504 31526 64518 31578
rect 64518 31526 64530 31578
rect 64530 31526 64560 31578
rect 64584 31526 64594 31578
rect 64594 31526 64640 31578
rect 64344 31524 64400 31526
rect 64424 31524 64480 31526
rect 64504 31524 64560 31526
rect 64584 31524 64640 31526
rect 64344 30490 64400 30492
rect 64424 30490 64480 30492
rect 64504 30490 64560 30492
rect 64584 30490 64640 30492
rect 64344 30438 64390 30490
rect 64390 30438 64400 30490
rect 64424 30438 64454 30490
rect 64454 30438 64466 30490
rect 64466 30438 64480 30490
rect 64504 30438 64518 30490
rect 64518 30438 64530 30490
rect 64530 30438 64560 30490
rect 64584 30438 64594 30490
rect 64594 30438 64640 30490
rect 64344 30436 64400 30438
rect 64424 30436 64480 30438
rect 64504 30436 64560 30438
rect 64584 30436 64640 30438
rect 64344 29402 64400 29404
rect 64424 29402 64480 29404
rect 64504 29402 64560 29404
rect 64584 29402 64640 29404
rect 64344 29350 64390 29402
rect 64390 29350 64400 29402
rect 64424 29350 64454 29402
rect 64454 29350 64466 29402
rect 64466 29350 64480 29402
rect 64504 29350 64518 29402
rect 64518 29350 64530 29402
rect 64530 29350 64560 29402
rect 64584 29350 64594 29402
rect 64594 29350 64640 29402
rect 64344 29348 64400 29350
rect 64424 29348 64480 29350
rect 64504 29348 64560 29350
rect 64584 29348 64640 29350
rect 65264 33210 65320 33212
rect 65344 33210 65400 33212
rect 65424 33210 65480 33212
rect 65504 33210 65560 33212
rect 65264 33158 65310 33210
rect 65310 33158 65320 33210
rect 65344 33158 65374 33210
rect 65374 33158 65386 33210
rect 65386 33158 65400 33210
rect 65424 33158 65438 33210
rect 65438 33158 65450 33210
rect 65450 33158 65480 33210
rect 65504 33158 65514 33210
rect 65514 33158 65560 33210
rect 65264 33156 65320 33158
rect 65344 33156 65400 33158
rect 65424 33156 65480 33158
rect 65504 33156 65560 33158
rect 65264 32122 65320 32124
rect 65344 32122 65400 32124
rect 65424 32122 65480 32124
rect 65504 32122 65560 32124
rect 65264 32070 65310 32122
rect 65310 32070 65320 32122
rect 65344 32070 65374 32122
rect 65374 32070 65386 32122
rect 65386 32070 65400 32122
rect 65424 32070 65438 32122
rect 65438 32070 65450 32122
rect 65450 32070 65480 32122
rect 65504 32070 65514 32122
rect 65514 32070 65560 32122
rect 65264 32068 65320 32070
rect 65344 32068 65400 32070
rect 65424 32068 65480 32070
rect 65504 32068 65560 32070
rect 64970 29008 65026 29064
rect 64878 28736 64934 28792
rect 64344 28314 64400 28316
rect 64424 28314 64480 28316
rect 64504 28314 64560 28316
rect 64584 28314 64640 28316
rect 64344 28262 64390 28314
rect 64390 28262 64400 28314
rect 64424 28262 64454 28314
rect 64454 28262 64466 28314
rect 64466 28262 64480 28314
rect 64504 28262 64518 28314
rect 64518 28262 64530 28314
rect 64530 28262 64560 28314
rect 64584 28262 64594 28314
rect 64594 28262 64640 28314
rect 64344 28260 64400 28262
rect 64424 28260 64480 28262
rect 64504 28260 64560 28262
rect 64584 28260 64640 28262
rect 64344 27226 64400 27228
rect 64424 27226 64480 27228
rect 64504 27226 64560 27228
rect 64584 27226 64640 27228
rect 64344 27174 64390 27226
rect 64390 27174 64400 27226
rect 64424 27174 64454 27226
rect 64454 27174 64466 27226
rect 64466 27174 64480 27226
rect 64504 27174 64518 27226
rect 64518 27174 64530 27226
rect 64530 27174 64560 27226
rect 64584 27174 64594 27226
rect 64594 27174 64640 27226
rect 64344 27172 64400 27174
rect 64424 27172 64480 27174
rect 64504 27172 64560 27174
rect 64584 27172 64640 27174
rect 64344 26138 64400 26140
rect 64424 26138 64480 26140
rect 64504 26138 64560 26140
rect 64584 26138 64640 26140
rect 64344 26086 64390 26138
rect 64390 26086 64400 26138
rect 64424 26086 64454 26138
rect 64454 26086 64466 26138
rect 64466 26086 64480 26138
rect 64504 26086 64518 26138
rect 64518 26086 64530 26138
rect 64530 26086 64560 26138
rect 64584 26086 64594 26138
rect 64594 26086 64640 26138
rect 64344 26084 64400 26086
rect 64424 26084 64480 26086
rect 64504 26084 64560 26086
rect 64584 26084 64640 26086
rect 64344 25050 64400 25052
rect 64424 25050 64480 25052
rect 64504 25050 64560 25052
rect 64584 25050 64640 25052
rect 64344 24998 64390 25050
rect 64390 24998 64400 25050
rect 64424 24998 64454 25050
rect 64454 24998 64466 25050
rect 64466 24998 64480 25050
rect 64504 24998 64518 25050
rect 64518 24998 64530 25050
rect 64530 24998 64560 25050
rect 64584 24998 64594 25050
rect 64594 24998 64640 25050
rect 64344 24996 64400 24998
rect 64424 24996 64480 24998
rect 64504 24996 64560 24998
rect 64584 24996 64640 24998
rect 65264 31034 65320 31036
rect 65344 31034 65400 31036
rect 65424 31034 65480 31036
rect 65504 31034 65560 31036
rect 65264 30982 65310 31034
rect 65310 30982 65320 31034
rect 65344 30982 65374 31034
rect 65374 30982 65386 31034
rect 65386 30982 65400 31034
rect 65424 30982 65438 31034
rect 65438 30982 65450 31034
rect 65450 30982 65480 31034
rect 65504 30982 65514 31034
rect 65514 30982 65560 31034
rect 65264 30980 65320 30982
rect 65344 30980 65400 30982
rect 65424 30980 65480 30982
rect 65504 30980 65560 30982
rect 66534 36624 66590 36680
rect 65264 29946 65320 29948
rect 65344 29946 65400 29948
rect 65424 29946 65480 29948
rect 65504 29946 65560 29948
rect 65264 29894 65310 29946
rect 65310 29894 65320 29946
rect 65344 29894 65374 29946
rect 65374 29894 65386 29946
rect 65386 29894 65400 29946
rect 65424 29894 65438 29946
rect 65438 29894 65450 29946
rect 65450 29894 65480 29946
rect 65504 29894 65514 29946
rect 65514 29894 65560 29946
rect 65264 29892 65320 29894
rect 65344 29892 65400 29894
rect 65424 29892 65480 29894
rect 65504 29892 65560 29894
rect 65264 28858 65320 28860
rect 65344 28858 65400 28860
rect 65424 28858 65480 28860
rect 65504 28858 65560 28860
rect 65264 28806 65310 28858
rect 65310 28806 65320 28858
rect 65344 28806 65374 28858
rect 65374 28806 65386 28858
rect 65386 28806 65400 28858
rect 65424 28806 65438 28858
rect 65438 28806 65450 28858
rect 65450 28806 65480 28858
rect 65504 28806 65514 28858
rect 65514 28806 65560 28858
rect 65264 28804 65320 28806
rect 65344 28804 65400 28806
rect 65424 28804 65480 28806
rect 65504 28804 65560 28806
rect 65264 27770 65320 27772
rect 65344 27770 65400 27772
rect 65424 27770 65480 27772
rect 65504 27770 65560 27772
rect 65264 27718 65310 27770
rect 65310 27718 65320 27770
rect 65344 27718 65374 27770
rect 65374 27718 65386 27770
rect 65386 27718 65400 27770
rect 65424 27718 65438 27770
rect 65438 27718 65450 27770
rect 65450 27718 65480 27770
rect 65504 27718 65514 27770
rect 65514 27718 65560 27770
rect 65264 27716 65320 27718
rect 65344 27716 65400 27718
rect 65424 27716 65480 27718
rect 65504 27716 65560 27718
rect 65264 26682 65320 26684
rect 65344 26682 65400 26684
rect 65424 26682 65480 26684
rect 65504 26682 65560 26684
rect 65264 26630 65310 26682
rect 65310 26630 65320 26682
rect 65344 26630 65374 26682
rect 65374 26630 65386 26682
rect 65386 26630 65400 26682
rect 65424 26630 65438 26682
rect 65438 26630 65450 26682
rect 65450 26630 65480 26682
rect 65504 26630 65514 26682
rect 65514 26630 65560 26682
rect 65264 26628 65320 26630
rect 65344 26628 65400 26630
rect 65424 26628 65480 26630
rect 65504 26628 65560 26630
rect 65264 25594 65320 25596
rect 65344 25594 65400 25596
rect 65424 25594 65480 25596
rect 65504 25594 65560 25596
rect 65264 25542 65310 25594
rect 65310 25542 65320 25594
rect 65344 25542 65374 25594
rect 65374 25542 65386 25594
rect 65386 25542 65400 25594
rect 65424 25542 65438 25594
rect 65438 25542 65450 25594
rect 65450 25542 65480 25594
rect 65504 25542 65514 25594
rect 65514 25542 65560 25594
rect 65264 25540 65320 25542
rect 65344 25540 65400 25542
rect 65424 25540 65480 25542
rect 65504 25540 65560 25542
rect 64344 23962 64400 23964
rect 64424 23962 64480 23964
rect 64504 23962 64560 23964
rect 64584 23962 64640 23964
rect 64344 23910 64390 23962
rect 64390 23910 64400 23962
rect 64424 23910 64454 23962
rect 64454 23910 64466 23962
rect 64466 23910 64480 23962
rect 64504 23910 64518 23962
rect 64518 23910 64530 23962
rect 64530 23910 64560 23962
rect 64584 23910 64594 23962
rect 64594 23910 64640 23962
rect 64344 23908 64400 23910
rect 64424 23908 64480 23910
rect 64504 23908 64560 23910
rect 64584 23908 64640 23910
rect 65264 24506 65320 24508
rect 65344 24506 65400 24508
rect 65424 24506 65480 24508
rect 65504 24506 65560 24508
rect 65264 24454 65310 24506
rect 65310 24454 65320 24506
rect 65344 24454 65374 24506
rect 65374 24454 65386 24506
rect 65386 24454 65400 24506
rect 65424 24454 65438 24506
rect 65438 24454 65450 24506
rect 65450 24454 65480 24506
rect 65504 24454 65514 24506
rect 65514 24454 65560 24506
rect 65264 24452 65320 24454
rect 65344 24452 65400 24454
rect 65424 24452 65480 24454
rect 65504 24452 65560 24454
rect 65264 23418 65320 23420
rect 65344 23418 65400 23420
rect 65424 23418 65480 23420
rect 65504 23418 65560 23420
rect 65264 23366 65310 23418
rect 65310 23366 65320 23418
rect 65344 23366 65374 23418
rect 65374 23366 65386 23418
rect 65386 23366 65400 23418
rect 65424 23366 65438 23418
rect 65438 23366 65450 23418
rect 65450 23366 65480 23418
rect 65504 23366 65514 23418
rect 65514 23366 65560 23418
rect 65264 23364 65320 23366
rect 65344 23364 65400 23366
rect 65424 23364 65480 23366
rect 65504 23364 65560 23366
rect 64344 22874 64400 22876
rect 64424 22874 64480 22876
rect 64504 22874 64560 22876
rect 64584 22874 64640 22876
rect 64344 22822 64390 22874
rect 64390 22822 64400 22874
rect 64424 22822 64454 22874
rect 64454 22822 64466 22874
rect 64466 22822 64480 22874
rect 64504 22822 64518 22874
rect 64518 22822 64530 22874
rect 64530 22822 64560 22874
rect 64584 22822 64594 22874
rect 64594 22822 64640 22874
rect 64344 22820 64400 22822
rect 64424 22820 64480 22822
rect 64504 22820 64560 22822
rect 64584 22820 64640 22822
rect 64344 21786 64400 21788
rect 64424 21786 64480 21788
rect 64504 21786 64560 21788
rect 64584 21786 64640 21788
rect 64344 21734 64390 21786
rect 64390 21734 64400 21786
rect 64424 21734 64454 21786
rect 64454 21734 64466 21786
rect 64466 21734 64480 21786
rect 64504 21734 64518 21786
rect 64518 21734 64530 21786
rect 64530 21734 64560 21786
rect 64584 21734 64594 21786
rect 64594 21734 64640 21786
rect 64344 21732 64400 21734
rect 64424 21732 64480 21734
rect 64504 21732 64560 21734
rect 64584 21732 64640 21734
rect 64344 20698 64400 20700
rect 64424 20698 64480 20700
rect 64504 20698 64560 20700
rect 64584 20698 64640 20700
rect 64344 20646 64390 20698
rect 64390 20646 64400 20698
rect 64424 20646 64454 20698
rect 64454 20646 64466 20698
rect 64466 20646 64480 20698
rect 64504 20646 64518 20698
rect 64518 20646 64530 20698
rect 64530 20646 64560 20698
rect 64584 20646 64594 20698
rect 64594 20646 64640 20698
rect 64344 20644 64400 20646
rect 64424 20644 64480 20646
rect 64504 20644 64560 20646
rect 64584 20644 64640 20646
rect 64344 19610 64400 19612
rect 64424 19610 64480 19612
rect 64504 19610 64560 19612
rect 64584 19610 64640 19612
rect 64344 19558 64390 19610
rect 64390 19558 64400 19610
rect 64424 19558 64454 19610
rect 64454 19558 64466 19610
rect 64466 19558 64480 19610
rect 64504 19558 64518 19610
rect 64518 19558 64530 19610
rect 64530 19558 64560 19610
rect 64584 19558 64594 19610
rect 64594 19558 64640 19610
rect 64344 19556 64400 19558
rect 64424 19556 64480 19558
rect 64504 19556 64560 19558
rect 64584 19556 64640 19558
rect 65264 22330 65320 22332
rect 65344 22330 65400 22332
rect 65424 22330 65480 22332
rect 65504 22330 65560 22332
rect 65264 22278 65310 22330
rect 65310 22278 65320 22330
rect 65344 22278 65374 22330
rect 65374 22278 65386 22330
rect 65386 22278 65400 22330
rect 65424 22278 65438 22330
rect 65438 22278 65450 22330
rect 65450 22278 65480 22330
rect 65504 22278 65514 22330
rect 65514 22278 65560 22330
rect 65264 22276 65320 22278
rect 65344 22276 65400 22278
rect 65424 22276 65480 22278
rect 65504 22276 65560 22278
rect 65264 21242 65320 21244
rect 65344 21242 65400 21244
rect 65424 21242 65480 21244
rect 65504 21242 65560 21244
rect 65264 21190 65310 21242
rect 65310 21190 65320 21242
rect 65344 21190 65374 21242
rect 65374 21190 65386 21242
rect 65386 21190 65400 21242
rect 65424 21190 65438 21242
rect 65438 21190 65450 21242
rect 65450 21190 65480 21242
rect 65504 21190 65514 21242
rect 65514 21190 65560 21242
rect 65264 21188 65320 21190
rect 65344 21188 65400 21190
rect 65424 21188 65480 21190
rect 65504 21188 65560 21190
rect 64344 18522 64400 18524
rect 64424 18522 64480 18524
rect 64504 18522 64560 18524
rect 64584 18522 64640 18524
rect 64344 18470 64390 18522
rect 64390 18470 64400 18522
rect 64424 18470 64454 18522
rect 64454 18470 64466 18522
rect 64466 18470 64480 18522
rect 64504 18470 64518 18522
rect 64518 18470 64530 18522
rect 64530 18470 64560 18522
rect 64584 18470 64594 18522
rect 64594 18470 64640 18522
rect 64344 18468 64400 18470
rect 64424 18468 64480 18470
rect 64504 18468 64560 18470
rect 64584 18468 64640 18470
rect 64344 17434 64400 17436
rect 64424 17434 64480 17436
rect 64504 17434 64560 17436
rect 64584 17434 64640 17436
rect 64344 17382 64390 17434
rect 64390 17382 64400 17434
rect 64424 17382 64454 17434
rect 64454 17382 64466 17434
rect 64466 17382 64480 17434
rect 64504 17382 64518 17434
rect 64518 17382 64530 17434
rect 64530 17382 64560 17434
rect 64584 17382 64594 17434
rect 64594 17382 64640 17434
rect 64344 17380 64400 17382
rect 64424 17380 64480 17382
rect 64504 17380 64560 17382
rect 64584 17380 64640 17382
rect 64344 16346 64400 16348
rect 64424 16346 64480 16348
rect 64504 16346 64560 16348
rect 64584 16346 64640 16348
rect 64344 16294 64390 16346
rect 64390 16294 64400 16346
rect 64424 16294 64454 16346
rect 64454 16294 64466 16346
rect 64466 16294 64480 16346
rect 64504 16294 64518 16346
rect 64518 16294 64530 16346
rect 64530 16294 64560 16346
rect 64584 16294 64594 16346
rect 64594 16294 64640 16346
rect 64344 16292 64400 16294
rect 64424 16292 64480 16294
rect 64504 16292 64560 16294
rect 64584 16292 64640 16294
rect 65264 20154 65320 20156
rect 65344 20154 65400 20156
rect 65424 20154 65480 20156
rect 65504 20154 65560 20156
rect 65264 20102 65310 20154
rect 65310 20102 65320 20154
rect 65344 20102 65374 20154
rect 65374 20102 65386 20154
rect 65386 20102 65400 20154
rect 65424 20102 65438 20154
rect 65438 20102 65450 20154
rect 65450 20102 65480 20154
rect 65504 20102 65514 20154
rect 65514 20102 65560 20154
rect 65264 20100 65320 20102
rect 65344 20100 65400 20102
rect 65424 20100 65480 20102
rect 65504 20100 65560 20102
rect 65264 19066 65320 19068
rect 65344 19066 65400 19068
rect 65424 19066 65480 19068
rect 65504 19066 65560 19068
rect 65264 19014 65310 19066
rect 65310 19014 65320 19066
rect 65344 19014 65374 19066
rect 65374 19014 65386 19066
rect 65386 19014 65400 19066
rect 65424 19014 65438 19066
rect 65438 19014 65450 19066
rect 65450 19014 65480 19066
rect 65504 19014 65514 19066
rect 65514 19014 65560 19066
rect 65264 19012 65320 19014
rect 65344 19012 65400 19014
rect 65424 19012 65480 19014
rect 65504 19012 65560 19014
rect 65264 17978 65320 17980
rect 65344 17978 65400 17980
rect 65424 17978 65480 17980
rect 65504 17978 65560 17980
rect 65264 17926 65310 17978
rect 65310 17926 65320 17978
rect 65344 17926 65374 17978
rect 65374 17926 65386 17978
rect 65386 17926 65400 17978
rect 65424 17926 65438 17978
rect 65438 17926 65450 17978
rect 65450 17926 65480 17978
rect 65504 17926 65514 17978
rect 65514 17926 65560 17978
rect 65264 17924 65320 17926
rect 65344 17924 65400 17926
rect 65424 17924 65480 17926
rect 65504 17924 65560 17926
rect 65264 16890 65320 16892
rect 65344 16890 65400 16892
rect 65424 16890 65480 16892
rect 65504 16890 65560 16892
rect 65264 16838 65310 16890
rect 65310 16838 65320 16890
rect 65344 16838 65374 16890
rect 65374 16838 65386 16890
rect 65386 16838 65400 16890
rect 65424 16838 65438 16890
rect 65438 16838 65450 16890
rect 65450 16838 65480 16890
rect 65504 16838 65514 16890
rect 65514 16838 65560 16890
rect 65264 16836 65320 16838
rect 65344 16836 65400 16838
rect 65424 16836 65480 16838
rect 65504 16836 65560 16838
rect 64970 16632 65026 16688
rect 64344 15258 64400 15260
rect 64424 15258 64480 15260
rect 64504 15258 64560 15260
rect 64584 15258 64640 15260
rect 64344 15206 64390 15258
rect 64390 15206 64400 15258
rect 64424 15206 64454 15258
rect 64454 15206 64466 15258
rect 64466 15206 64480 15258
rect 64504 15206 64518 15258
rect 64518 15206 64530 15258
rect 64530 15206 64560 15258
rect 64584 15206 64594 15258
rect 64594 15206 64640 15258
rect 64344 15204 64400 15206
rect 64424 15204 64480 15206
rect 64504 15204 64560 15206
rect 64584 15204 64640 15206
rect 64142 15136 64198 15192
rect 64344 14170 64400 14172
rect 64424 14170 64480 14172
rect 64504 14170 64560 14172
rect 64584 14170 64640 14172
rect 64344 14118 64390 14170
rect 64390 14118 64400 14170
rect 64424 14118 64454 14170
rect 64454 14118 64466 14170
rect 64466 14118 64480 14170
rect 64504 14118 64518 14170
rect 64518 14118 64530 14170
rect 64530 14118 64560 14170
rect 64584 14118 64594 14170
rect 64594 14118 64640 14170
rect 64344 14116 64400 14118
rect 64424 14116 64480 14118
rect 64504 14116 64560 14118
rect 64584 14116 64640 14118
rect 64344 13082 64400 13084
rect 64424 13082 64480 13084
rect 64504 13082 64560 13084
rect 64584 13082 64640 13084
rect 64344 13030 64390 13082
rect 64390 13030 64400 13082
rect 64424 13030 64454 13082
rect 64454 13030 64466 13082
rect 64466 13030 64480 13082
rect 64504 13030 64518 13082
rect 64518 13030 64530 13082
rect 64530 13030 64560 13082
rect 64584 13030 64594 13082
rect 64594 13030 64640 13082
rect 64344 13028 64400 13030
rect 64424 13028 64480 13030
rect 64504 13028 64560 13030
rect 64584 13028 64640 13030
rect 64344 11994 64400 11996
rect 64424 11994 64480 11996
rect 64504 11994 64560 11996
rect 64584 11994 64640 11996
rect 64344 11942 64390 11994
rect 64390 11942 64400 11994
rect 64424 11942 64454 11994
rect 64454 11942 64466 11994
rect 64466 11942 64480 11994
rect 64504 11942 64518 11994
rect 64518 11942 64530 11994
rect 64530 11942 64560 11994
rect 64584 11942 64594 11994
rect 64594 11942 64640 11994
rect 64344 11940 64400 11942
rect 64424 11940 64480 11942
rect 64504 11940 64560 11942
rect 64584 11940 64640 11942
rect 64344 10906 64400 10908
rect 64424 10906 64480 10908
rect 64504 10906 64560 10908
rect 64584 10906 64640 10908
rect 64344 10854 64390 10906
rect 64390 10854 64400 10906
rect 64424 10854 64454 10906
rect 64454 10854 64466 10906
rect 64466 10854 64480 10906
rect 64504 10854 64518 10906
rect 64518 10854 64530 10906
rect 64530 10854 64560 10906
rect 64584 10854 64594 10906
rect 64594 10854 64640 10906
rect 64344 10852 64400 10854
rect 64424 10852 64480 10854
rect 64504 10852 64560 10854
rect 64584 10852 64640 10854
rect 64344 9818 64400 9820
rect 64424 9818 64480 9820
rect 64504 9818 64560 9820
rect 64584 9818 64640 9820
rect 64344 9766 64390 9818
rect 64390 9766 64400 9818
rect 64424 9766 64454 9818
rect 64454 9766 64466 9818
rect 64466 9766 64480 9818
rect 64504 9766 64518 9818
rect 64518 9766 64530 9818
rect 64530 9766 64560 9818
rect 64584 9766 64594 9818
rect 64594 9766 64640 9818
rect 64344 9764 64400 9766
rect 64424 9764 64480 9766
rect 64504 9764 64560 9766
rect 64584 9764 64640 9766
rect 64344 8730 64400 8732
rect 64424 8730 64480 8732
rect 64504 8730 64560 8732
rect 64584 8730 64640 8732
rect 64344 8678 64390 8730
rect 64390 8678 64400 8730
rect 64424 8678 64454 8730
rect 64454 8678 64466 8730
rect 64466 8678 64480 8730
rect 64504 8678 64518 8730
rect 64518 8678 64530 8730
rect 64530 8678 64560 8730
rect 64584 8678 64594 8730
rect 64594 8678 64640 8730
rect 64344 8676 64400 8678
rect 64424 8676 64480 8678
rect 64504 8676 64560 8678
rect 64584 8676 64640 8678
rect 64344 7642 64400 7644
rect 64424 7642 64480 7644
rect 64504 7642 64560 7644
rect 64584 7642 64640 7644
rect 64344 7590 64390 7642
rect 64390 7590 64400 7642
rect 64424 7590 64454 7642
rect 64454 7590 64466 7642
rect 64466 7590 64480 7642
rect 64504 7590 64518 7642
rect 64518 7590 64530 7642
rect 64530 7590 64560 7642
rect 64584 7590 64594 7642
rect 64594 7590 64640 7642
rect 64344 7588 64400 7590
rect 64424 7588 64480 7590
rect 64504 7588 64560 7590
rect 64584 7588 64640 7590
rect 65264 15802 65320 15804
rect 65344 15802 65400 15804
rect 65424 15802 65480 15804
rect 65504 15802 65560 15804
rect 65264 15750 65310 15802
rect 65310 15750 65320 15802
rect 65344 15750 65374 15802
rect 65374 15750 65386 15802
rect 65386 15750 65400 15802
rect 65424 15750 65438 15802
rect 65438 15750 65450 15802
rect 65450 15750 65480 15802
rect 65504 15750 65514 15802
rect 65514 15750 65560 15802
rect 65264 15748 65320 15750
rect 65344 15748 65400 15750
rect 65424 15748 65480 15750
rect 65504 15748 65560 15750
rect 65264 14714 65320 14716
rect 65344 14714 65400 14716
rect 65424 14714 65480 14716
rect 65504 14714 65560 14716
rect 65264 14662 65310 14714
rect 65310 14662 65320 14714
rect 65344 14662 65374 14714
rect 65374 14662 65386 14714
rect 65386 14662 65400 14714
rect 65424 14662 65438 14714
rect 65438 14662 65450 14714
rect 65450 14662 65480 14714
rect 65504 14662 65514 14714
rect 65514 14662 65560 14714
rect 65264 14660 65320 14662
rect 65344 14660 65400 14662
rect 65424 14660 65480 14662
rect 65504 14660 65560 14662
rect 65264 13626 65320 13628
rect 65344 13626 65400 13628
rect 65424 13626 65480 13628
rect 65504 13626 65560 13628
rect 65264 13574 65310 13626
rect 65310 13574 65320 13626
rect 65344 13574 65374 13626
rect 65374 13574 65386 13626
rect 65386 13574 65400 13626
rect 65424 13574 65438 13626
rect 65438 13574 65450 13626
rect 65450 13574 65480 13626
rect 65504 13574 65514 13626
rect 65514 13574 65560 13626
rect 65264 13572 65320 13574
rect 65344 13572 65400 13574
rect 65424 13572 65480 13574
rect 65504 13572 65560 13574
rect 66074 16632 66130 16688
rect 65264 12538 65320 12540
rect 65344 12538 65400 12540
rect 65424 12538 65480 12540
rect 65504 12538 65560 12540
rect 65264 12486 65310 12538
rect 65310 12486 65320 12538
rect 65344 12486 65374 12538
rect 65374 12486 65386 12538
rect 65386 12486 65400 12538
rect 65424 12486 65438 12538
rect 65438 12486 65450 12538
rect 65450 12486 65480 12538
rect 65504 12486 65514 12538
rect 65514 12486 65560 12538
rect 65264 12484 65320 12486
rect 65344 12484 65400 12486
rect 65424 12484 65480 12486
rect 65504 12484 65560 12486
rect 65264 11450 65320 11452
rect 65344 11450 65400 11452
rect 65424 11450 65480 11452
rect 65504 11450 65560 11452
rect 65264 11398 65310 11450
rect 65310 11398 65320 11450
rect 65344 11398 65374 11450
rect 65374 11398 65386 11450
rect 65386 11398 65400 11450
rect 65424 11398 65438 11450
rect 65438 11398 65450 11450
rect 65450 11398 65480 11450
rect 65504 11398 65514 11450
rect 65514 11398 65560 11450
rect 65264 11396 65320 11398
rect 65344 11396 65400 11398
rect 65424 11396 65480 11398
rect 65504 11396 65560 11398
rect 65264 10362 65320 10364
rect 65344 10362 65400 10364
rect 65424 10362 65480 10364
rect 65504 10362 65560 10364
rect 65264 10310 65310 10362
rect 65310 10310 65320 10362
rect 65344 10310 65374 10362
rect 65374 10310 65386 10362
rect 65386 10310 65400 10362
rect 65424 10310 65438 10362
rect 65438 10310 65450 10362
rect 65450 10310 65480 10362
rect 65504 10310 65514 10362
rect 65514 10310 65560 10362
rect 65264 10308 65320 10310
rect 65344 10308 65400 10310
rect 65424 10308 65480 10310
rect 65504 10308 65560 10310
rect 65264 9274 65320 9276
rect 65344 9274 65400 9276
rect 65424 9274 65480 9276
rect 65504 9274 65560 9276
rect 65264 9222 65310 9274
rect 65310 9222 65320 9274
rect 65344 9222 65374 9274
rect 65374 9222 65386 9274
rect 65386 9222 65400 9274
rect 65424 9222 65438 9274
rect 65438 9222 65450 9274
rect 65450 9222 65480 9274
rect 65504 9222 65514 9274
rect 65514 9222 65560 9274
rect 65264 9220 65320 9222
rect 65344 9220 65400 9222
rect 65424 9220 65480 9222
rect 65504 9220 65560 9222
rect 64142 5908 64198 5944
rect 64142 5888 64144 5908
rect 64144 5888 64196 5908
rect 64196 5888 64198 5908
rect 64344 6554 64400 6556
rect 64424 6554 64480 6556
rect 64504 6554 64560 6556
rect 64584 6554 64640 6556
rect 64344 6502 64390 6554
rect 64390 6502 64400 6554
rect 64424 6502 64454 6554
rect 64454 6502 64466 6554
rect 64466 6502 64480 6554
rect 64504 6502 64518 6554
rect 64518 6502 64530 6554
rect 64530 6502 64560 6554
rect 64584 6502 64594 6554
rect 64594 6502 64640 6554
rect 64344 6500 64400 6502
rect 64424 6500 64480 6502
rect 64504 6500 64560 6502
rect 64584 6500 64640 6502
rect 64694 6060 64696 6080
rect 64696 6060 64748 6080
rect 64748 6060 64750 6080
rect 64694 6024 64750 6060
rect 64344 5466 64400 5468
rect 64424 5466 64480 5468
rect 64504 5466 64560 5468
rect 64584 5466 64640 5468
rect 64344 5414 64390 5466
rect 64390 5414 64400 5466
rect 64424 5414 64454 5466
rect 64454 5414 64466 5466
rect 64466 5414 64480 5466
rect 64504 5414 64518 5466
rect 64518 5414 64530 5466
rect 64530 5414 64560 5466
rect 64584 5414 64594 5466
rect 64594 5414 64640 5466
rect 64344 5412 64400 5414
rect 64424 5412 64480 5414
rect 64504 5412 64560 5414
rect 64584 5412 64640 5414
rect 64344 4378 64400 4380
rect 64424 4378 64480 4380
rect 64504 4378 64560 4380
rect 64584 4378 64640 4380
rect 64344 4326 64390 4378
rect 64390 4326 64400 4378
rect 64424 4326 64454 4378
rect 64454 4326 64466 4378
rect 64466 4326 64480 4378
rect 64504 4326 64518 4378
rect 64518 4326 64530 4378
rect 64530 4326 64560 4378
rect 64584 4326 64594 4378
rect 64594 4326 64640 4378
rect 64344 4324 64400 4326
rect 64424 4324 64480 4326
rect 64504 4324 64560 4326
rect 64584 4324 64640 4326
rect 64344 3290 64400 3292
rect 64424 3290 64480 3292
rect 64504 3290 64560 3292
rect 64584 3290 64640 3292
rect 64344 3238 64390 3290
rect 64390 3238 64400 3290
rect 64424 3238 64454 3290
rect 64454 3238 64466 3290
rect 64466 3238 64480 3290
rect 64504 3238 64518 3290
rect 64518 3238 64530 3290
rect 64530 3238 64560 3290
rect 64584 3238 64594 3290
rect 64594 3238 64640 3290
rect 64344 3236 64400 3238
rect 64424 3236 64480 3238
rect 64504 3236 64560 3238
rect 64584 3236 64640 3238
rect 64344 2202 64400 2204
rect 64424 2202 64480 2204
rect 64504 2202 64560 2204
rect 64584 2202 64640 2204
rect 64344 2150 64390 2202
rect 64390 2150 64400 2202
rect 64424 2150 64454 2202
rect 64454 2150 64466 2202
rect 64466 2150 64480 2202
rect 64504 2150 64518 2202
rect 64518 2150 64530 2202
rect 64530 2150 64560 2202
rect 64584 2150 64594 2202
rect 64594 2150 64640 2202
rect 64344 2148 64400 2150
rect 64424 2148 64480 2150
rect 64504 2148 64560 2150
rect 64584 2148 64640 2150
rect 64694 1944 64750 2000
rect 63498 1808 63554 1864
rect 62854 1536 62910 1592
rect 62578 1264 62634 1320
rect 64344 1114 64400 1116
rect 64424 1114 64480 1116
rect 64504 1114 64560 1116
rect 64584 1114 64640 1116
rect 64344 1062 64390 1114
rect 64390 1062 64400 1114
rect 64424 1062 64454 1114
rect 64454 1062 64466 1114
rect 64466 1062 64480 1114
rect 64504 1062 64518 1114
rect 64518 1062 64530 1114
rect 64530 1062 64560 1114
rect 64584 1062 64594 1114
rect 64594 1062 64640 1114
rect 64344 1060 64400 1062
rect 64424 1060 64480 1062
rect 64504 1060 64560 1062
rect 64584 1060 64640 1062
rect 65264 8186 65320 8188
rect 65344 8186 65400 8188
rect 65424 8186 65480 8188
rect 65504 8186 65560 8188
rect 65264 8134 65310 8186
rect 65310 8134 65320 8186
rect 65344 8134 65374 8186
rect 65374 8134 65386 8186
rect 65386 8134 65400 8186
rect 65424 8134 65438 8186
rect 65438 8134 65450 8186
rect 65450 8134 65480 8186
rect 65504 8134 65514 8186
rect 65514 8134 65560 8186
rect 65264 8132 65320 8134
rect 65344 8132 65400 8134
rect 65424 8132 65480 8134
rect 65504 8132 65560 8134
rect 65264 7098 65320 7100
rect 65344 7098 65400 7100
rect 65424 7098 65480 7100
rect 65504 7098 65560 7100
rect 65264 7046 65310 7098
rect 65310 7046 65320 7098
rect 65344 7046 65374 7098
rect 65374 7046 65386 7098
rect 65386 7046 65400 7098
rect 65424 7046 65438 7098
rect 65438 7046 65450 7098
rect 65450 7046 65480 7098
rect 65504 7046 65514 7098
rect 65514 7046 65560 7098
rect 65264 7044 65320 7046
rect 65344 7044 65400 7046
rect 65424 7044 65480 7046
rect 65504 7044 65560 7046
rect 65264 6010 65320 6012
rect 65344 6010 65400 6012
rect 65424 6010 65480 6012
rect 65504 6010 65560 6012
rect 65264 5958 65310 6010
rect 65310 5958 65320 6010
rect 65344 5958 65374 6010
rect 65374 5958 65386 6010
rect 65386 5958 65400 6010
rect 65424 5958 65438 6010
rect 65438 5958 65450 6010
rect 65450 5958 65480 6010
rect 65504 5958 65514 6010
rect 65514 5958 65560 6010
rect 65264 5956 65320 5958
rect 65344 5956 65400 5958
rect 65424 5956 65480 5958
rect 65504 5956 65560 5958
rect 65264 4922 65320 4924
rect 65344 4922 65400 4924
rect 65424 4922 65480 4924
rect 65504 4922 65560 4924
rect 65264 4870 65310 4922
rect 65310 4870 65320 4922
rect 65344 4870 65374 4922
rect 65374 4870 65386 4922
rect 65386 4870 65400 4922
rect 65424 4870 65438 4922
rect 65438 4870 65450 4922
rect 65450 4870 65480 4922
rect 65504 4870 65514 4922
rect 65514 4870 65560 4922
rect 65264 4868 65320 4870
rect 65344 4868 65400 4870
rect 65424 4868 65480 4870
rect 65504 4868 65560 4870
rect 65264 3834 65320 3836
rect 65344 3834 65400 3836
rect 65424 3834 65480 3836
rect 65504 3834 65560 3836
rect 65264 3782 65310 3834
rect 65310 3782 65320 3834
rect 65344 3782 65374 3834
rect 65374 3782 65386 3834
rect 65386 3782 65400 3834
rect 65424 3782 65438 3834
rect 65438 3782 65450 3834
rect 65450 3782 65480 3834
rect 65504 3782 65514 3834
rect 65514 3782 65560 3834
rect 65264 3780 65320 3782
rect 65344 3780 65400 3782
rect 65424 3780 65480 3782
rect 65504 3780 65560 3782
rect 65264 2746 65320 2748
rect 65344 2746 65400 2748
rect 65424 2746 65480 2748
rect 65504 2746 65560 2748
rect 65264 2694 65310 2746
rect 65310 2694 65320 2746
rect 65344 2694 65374 2746
rect 65374 2694 65386 2746
rect 65386 2694 65400 2746
rect 65424 2694 65438 2746
rect 65438 2694 65450 2746
rect 65450 2694 65480 2746
rect 65504 2694 65514 2746
rect 65514 2694 65560 2746
rect 65264 2692 65320 2694
rect 65344 2692 65400 2694
rect 65424 2692 65480 2694
rect 65504 2692 65560 2694
rect 65264 1658 65320 1660
rect 65344 1658 65400 1660
rect 65424 1658 65480 1660
rect 65504 1658 65560 1660
rect 65264 1606 65310 1658
rect 65310 1606 65320 1658
rect 65344 1606 65374 1658
rect 65374 1606 65386 1658
rect 65386 1606 65400 1658
rect 65424 1606 65438 1658
rect 65438 1606 65450 1658
rect 65450 1606 65480 1658
rect 65504 1606 65514 1658
rect 65514 1606 65560 1658
rect 65264 1604 65320 1606
rect 65344 1604 65400 1606
rect 65424 1604 65480 1606
rect 65504 1604 65560 1606
rect 65264 570 65320 572
rect 65344 570 65400 572
rect 65424 570 65480 572
rect 65504 570 65560 572
rect 65264 518 65310 570
rect 65310 518 65320 570
rect 65344 518 65374 570
rect 65374 518 65386 570
rect 65386 518 65400 570
rect 65424 518 65438 570
rect 65438 518 65450 570
rect 65450 518 65480 570
rect 65504 518 65514 570
rect 65514 518 65560 570
rect 65264 516 65320 518
rect 65344 516 65400 518
rect 65424 516 65480 518
rect 65504 516 65560 518
<< metal3 >>
rect 35341 45114 35407 45117
rect 26006 45112 35407 45114
rect 26006 45056 35346 45112
rect 35402 45056 35407 45112
rect 26006 45054 35407 45056
rect 24342 44916 24348 44980
rect 24412 44978 24418 44980
rect 24853 44978 24919 44981
rect 26006 44980 26066 45054
rect 35341 45051 35407 45054
rect 24412 44976 24919 44978
rect 24412 44920 24858 44976
rect 24914 44920 24919 44976
rect 24412 44918 24919 44920
rect 24412 44916 24418 44918
rect 24853 44915 24919 44918
rect 25998 44916 26004 44980
rect 26068 44916 26074 44980
rect 25446 44780 25452 44844
rect 25516 44842 25522 44844
rect 31753 44842 31819 44845
rect 25516 44840 31819 44842
rect 25516 44784 31758 44840
rect 31814 44784 31819 44840
rect 25516 44782 31819 44784
rect 25516 44780 25522 44782
rect 31753 44779 31819 44782
rect 11646 44644 11652 44708
rect 11716 44706 11722 44708
rect 12525 44706 12591 44709
rect 11716 44704 12591 44706
rect 11716 44648 12530 44704
rect 12586 44648 12591 44704
rect 11716 44646 12591 44648
rect 11716 44644 11722 44646
rect 12525 44643 12591 44646
rect 14958 44644 14964 44708
rect 15028 44706 15034 44708
rect 16205 44706 16271 44709
rect 15028 44704 16271 44706
rect 15028 44648 16210 44704
rect 16266 44648 16271 44704
rect 15028 44646 16271 44648
rect 15028 44644 15034 44646
rect 16205 44643 16271 44646
rect 17217 44706 17283 44709
rect 17718 44706 17724 44708
rect 17217 44704 17724 44706
rect 17217 44648 17222 44704
rect 17278 44648 17724 44704
rect 17217 44646 17724 44648
rect 17217 44643 17283 44646
rect 17718 44644 17724 44646
rect 17788 44644 17794 44708
rect 26601 44706 26667 44709
rect 27654 44706 27660 44708
rect 26601 44704 27660 44706
rect 26601 44648 26606 44704
rect 26662 44648 27660 44704
rect 26601 44646 27660 44648
rect 26601 44643 26667 44646
rect 27654 44644 27660 44646
rect 27724 44644 27730 44708
rect 1994 44640 2310 44641
rect 1994 44576 2000 44640
rect 2064 44576 2080 44640
rect 2144 44576 2160 44640
rect 2224 44576 2240 44640
rect 2304 44576 2310 44640
rect 1994 44575 2310 44576
rect 50994 44640 51310 44641
rect 50994 44576 51000 44640
rect 51064 44576 51080 44640
rect 51144 44576 51160 44640
rect 51224 44576 51240 44640
rect 51304 44576 51310 44640
rect 50994 44575 51310 44576
rect 6177 44572 6243 44573
rect 6729 44572 6795 44573
rect 7281 44572 7347 44573
rect 7833 44572 7899 44573
rect 8385 44572 8451 44573
rect 8937 44572 9003 44573
rect 9489 44572 9555 44573
rect 10041 44572 10107 44573
rect 10593 44572 10659 44573
rect 12249 44572 12315 44573
rect 12801 44572 12867 44573
rect 6126 44508 6132 44572
rect 6196 44570 6243 44572
rect 6196 44568 6288 44570
rect 6238 44512 6288 44568
rect 6196 44510 6288 44512
rect 6196 44508 6243 44510
rect 6678 44508 6684 44572
rect 6748 44570 6795 44572
rect 6748 44568 6840 44570
rect 6790 44512 6840 44568
rect 6748 44510 6840 44512
rect 6748 44508 6795 44510
rect 7230 44508 7236 44572
rect 7300 44570 7347 44572
rect 7300 44568 7392 44570
rect 7342 44512 7392 44568
rect 7300 44510 7392 44512
rect 7300 44508 7347 44510
rect 7782 44508 7788 44572
rect 7852 44570 7899 44572
rect 7852 44568 7944 44570
rect 7894 44512 7944 44568
rect 7852 44510 7944 44512
rect 7852 44508 7899 44510
rect 8334 44508 8340 44572
rect 8404 44570 8451 44572
rect 8404 44568 8496 44570
rect 8446 44512 8496 44568
rect 8404 44510 8496 44512
rect 8404 44508 8451 44510
rect 8886 44508 8892 44572
rect 8956 44570 9003 44572
rect 8956 44568 9048 44570
rect 8998 44512 9048 44568
rect 8956 44510 9048 44512
rect 8956 44508 9003 44510
rect 9438 44508 9444 44572
rect 9508 44570 9555 44572
rect 9508 44568 9600 44570
rect 9550 44512 9600 44568
rect 9508 44510 9600 44512
rect 9508 44508 9555 44510
rect 9990 44508 9996 44572
rect 10060 44570 10107 44572
rect 10060 44568 10152 44570
rect 10102 44512 10152 44568
rect 10060 44510 10152 44512
rect 10060 44508 10107 44510
rect 10542 44508 10548 44572
rect 10612 44570 10659 44572
rect 10612 44568 10704 44570
rect 10654 44512 10704 44568
rect 10612 44510 10704 44512
rect 10612 44508 10659 44510
rect 12198 44508 12204 44572
rect 12268 44570 12315 44572
rect 12268 44568 12360 44570
rect 12310 44512 12360 44568
rect 12268 44510 12360 44512
rect 12268 44508 12315 44510
rect 12750 44508 12756 44572
rect 12820 44570 12867 44572
rect 12820 44568 12912 44570
rect 12862 44512 12912 44568
rect 12820 44510 12912 44512
rect 12820 44508 12867 44510
rect 13302 44508 13308 44572
rect 13372 44570 13378 44572
rect 13537 44570 13603 44573
rect 13813 44572 13879 44573
rect 15469 44572 15535 44573
rect 13813 44570 13860 44572
rect 13372 44568 13603 44570
rect 13372 44512 13542 44568
rect 13598 44512 13603 44568
rect 13372 44510 13603 44512
rect 13768 44568 13860 44570
rect 13768 44512 13818 44568
rect 13768 44510 13860 44512
rect 13372 44508 13378 44510
rect 6177 44507 6243 44508
rect 6729 44507 6795 44508
rect 7281 44507 7347 44508
rect 7833 44507 7899 44508
rect 8385 44507 8451 44508
rect 8937 44507 9003 44508
rect 9489 44507 9555 44508
rect 10041 44507 10107 44508
rect 10593 44507 10659 44508
rect 12249 44507 12315 44508
rect 12801 44507 12867 44508
rect 13537 44507 13603 44510
rect 13813 44508 13860 44510
rect 13924 44508 13930 44572
rect 15469 44570 15516 44572
rect 15424 44568 15516 44570
rect 15424 44512 15474 44568
rect 15424 44510 15516 44512
rect 15469 44508 15516 44510
rect 15580 44508 15586 44572
rect 15929 44570 15995 44573
rect 16665 44572 16731 44573
rect 16062 44570 16068 44572
rect 15929 44568 16068 44570
rect 15929 44512 15934 44568
rect 15990 44512 16068 44568
rect 15929 44510 16068 44512
rect 13813 44507 13879 44508
rect 15469 44507 15535 44508
rect 15929 44507 15995 44510
rect 16062 44508 16068 44510
rect 16132 44508 16138 44572
rect 16614 44508 16620 44572
rect 16684 44570 16731 44572
rect 16941 44570 17007 44573
rect 17166 44570 17172 44572
rect 16684 44568 16776 44570
rect 16726 44512 16776 44568
rect 16684 44510 16776 44512
rect 16941 44568 17172 44570
rect 16941 44512 16946 44568
rect 17002 44512 17172 44568
rect 16941 44510 17172 44512
rect 16684 44508 16731 44510
rect 16665 44507 16731 44508
rect 16941 44507 17007 44510
rect 17166 44508 17172 44510
rect 17236 44508 17242 44572
rect 26233 44434 26299 44437
rect 26550 44434 26556 44436
rect 26233 44432 26556 44434
rect 26233 44376 26238 44432
rect 26294 44376 26556 44432
rect 26233 44374 26556 44376
rect 26233 44371 26299 44374
rect 26550 44372 26556 44374
rect 26620 44372 26626 44436
rect 26785 44434 26851 44437
rect 27102 44434 27108 44436
rect 26785 44432 27108 44434
rect 26785 44376 26790 44432
rect 26846 44376 27108 44432
rect 26785 44374 27108 44376
rect 26785 44371 26851 44374
rect 27102 44372 27108 44374
rect 27172 44372 27178 44436
rect 27521 44434 27587 44437
rect 28206 44434 28212 44436
rect 27521 44432 28212 44434
rect 27521 44376 27526 44432
rect 27582 44376 28212 44432
rect 27521 44374 28212 44376
rect 27521 44371 27587 44374
rect 28206 44372 28212 44374
rect 28276 44372 28282 44436
rect 2914 44096 3230 44097
rect 2914 44032 2920 44096
rect 2984 44032 3000 44096
rect 3064 44032 3080 44096
rect 3144 44032 3160 44096
rect 3224 44032 3230 44096
rect 2914 44031 3230 44032
rect 51914 44096 52230 44097
rect 51914 44032 51920 44096
rect 51984 44032 52000 44096
rect 52064 44032 52080 44096
rect 52144 44032 52160 44096
rect 52224 44032 52230 44096
rect 51914 44031 52230 44032
rect 11145 43892 11211 43893
rect 11094 43828 11100 43892
rect 11164 43890 11211 43892
rect 11164 43888 11256 43890
rect 11206 43832 11256 43888
rect 11164 43830 11256 43832
rect 11164 43828 11211 43830
rect 14406 43828 14412 43892
rect 14476 43890 14482 43892
rect 15285 43890 15351 43893
rect 14476 43888 15351 43890
rect 14476 43832 15290 43888
rect 15346 43832 15351 43888
rect 14476 43830 15351 43832
rect 14476 43828 14482 43830
rect 11145 43827 11211 43828
rect 15285 43827 15351 43830
rect 17953 43754 18019 43757
rect 18822 43754 18828 43756
rect 17953 43752 18828 43754
rect 17953 43696 17958 43752
rect 18014 43696 18828 43752
rect 17953 43694 18828 43696
rect 17953 43691 18019 43694
rect 18822 43692 18828 43694
rect 18892 43692 18898 43756
rect 19793 43754 19859 43757
rect 26509 43754 26575 43757
rect 19793 43752 26575 43754
rect 19793 43696 19798 43752
rect 19854 43696 26514 43752
rect 26570 43696 26575 43752
rect 19793 43694 26575 43696
rect 19793 43691 19859 43694
rect 26509 43691 26575 43694
rect 31385 43754 31451 43757
rect 31886 43754 31892 43756
rect 31385 43752 31892 43754
rect 31385 43696 31390 43752
rect 31446 43696 31892 43752
rect 31385 43694 31892 43696
rect 31385 43691 31451 43694
rect 31886 43692 31892 43694
rect 31956 43692 31962 43756
rect 1994 43552 2310 43553
rect 1994 43488 2000 43552
rect 2064 43488 2080 43552
rect 2144 43488 2160 43552
rect 2224 43488 2240 43552
rect 2304 43488 2310 43552
rect 1994 43487 2310 43488
rect 50994 43552 51310 43553
rect 50994 43488 51000 43552
rect 51064 43488 51080 43552
rect 51144 43488 51160 43552
rect 51224 43488 51240 43552
rect 51304 43488 51310 43552
rect 50994 43487 51310 43488
rect 18270 43420 18276 43484
rect 18340 43482 18346 43484
rect 18781 43482 18847 43485
rect 18340 43480 18847 43482
rect 18340 43424 18786 43480
rect 18842 43424 18847 43480
rect 18340 43422 18847 43424
rect 18340 43420 18346 43422
rect 18781 43419 18847 43422
rect 30557 43482 30623 43485
rect 31661 43482 31727 43485
rect 30557 43480 31727 43482
rect 30557 43424 30562 43480
rect 30618 43424 31666 43480
rect 31722 43424 31727 43480
rect 30557 43422 31727 43424
rect 30557 43419 30623 43422
rect 31661 43419 31727 43422
rect 29637 43346 29703 43349
rect 31201 43346 31267 43349
rect 29637 43344 31267 43346
rect 29637 43288 29642 43344
rect 29698 43288 31206 43344
rect 31262 43288 31267 43344
rect 29637 43286 31267 43288
rect 29637 43283 29703 43286
rect 31201 43283 31267 43286
rect 22686 43148 22692 43212
rect 22756 43210 22762 43212
rect 24526 43210 24532 43212
rect 22756 43150 24532 43210
rect 22756 43148 22762 43150
rect 24526 43148 24532 43150
rect 24596 43148 24602 43212
rect 27102 43012 27108 43076
rect 27172 43074 27178 43076
rect 36813 43074 36879 43077
rect 27172 43072 36879 43074
rect 27172 43016 36818 43072
rect 36874 43016 36879 43072
rect 27172 43014 36879 43016
rect 27172 43012 27178 43014
rect 36813 43011 36879 43014
rect 2914 43008 3230 43009
rect 2914 42944 2920 43008
rect 2984 42944 3000 43008
rect 3064 42944 3080 43008
rect 3144 42944 3160 43008
rect 3224 42944 3230 43008
rect 2914 42943 3230 42944
rect 51914 43008 52230 43009
rect 51914 42944 51920 43008
rect 51984 42944 52000 43008
rect 52064 42944 52080 43008
rect 52144 42944 52160 43008
rect 52224 42944 52230 43008
rect 51914 42943 52230 42944
rect 23238 42740 23244 42804
rect 23308 42802 23314 42804
rect 28942 42802 28948 42804
rect 23308 42742 28948 42802
rect 23308 42740 23314 42742
rect 28942 42740 28948 42742
rect 29012 42740 29018 42804
rect 26601 42666 26667 42669
rect 27797 42666 27863 42669
rect 26601 42664 27863 42666
rect 26601 42608 26606 42664
rect 26662 42608 27802 42664
rect 27858 42608 27863 42664
rect 26601 42606 27863 42608
rect 26601 42603 26667 42606
rect 27797 42603 27863 42606
rect 31845 42666 31911 42669
rect 60733 42666 60799 42669
rect 31845 42664 60799 42666
rect 31845 42608 31850 42664
rect 31906 42608 60738 42664
rect 60794 42608 60799 42664
rect 31845 42606 60799 42608
rect 31845 42603 31911 42606
rect 60733 42603 60799 42606
rect 32489 42530 32555 42533
rect 22050 42528 32555 42530
rect 22050 42472 32494 42528
rect 32550 42472 32555 42528
rect 22050 42470 32555 42472
rect 1994 42464 2310 42465
rect 1994 42400 2000 42464
rect 2064 42400 2080 42464
rect 2144 42400 2160 42464
rect 2224 42400 2240 42464
rect 2304 42400 2310 42464
rect 1994 42399 2310 42400
rect 16849 42258 16915 42261
rect 22050 42258 22110 42470
rect 32489 42467 32555 42470
rect 50994 42464 51310 42465
rect 50994 42400 51000 42464
rect 51064 42400 51080 42464
rect 51144 42400 51160 42464
rect 51224 42400 51240 42464
rect 51304 42400 51310 42464
rect 50994 42399 51310 42400
rect 27838 42332 27844 42396
rect 27908 42394 27914 42396
rect 35065 42394 35131 42397
rect 27908 42392 35131 42394
rect 27908 42336 35070 42392
rect 35126 42336 35131 42392
rect 27908 42334 35131 42336
rect 27908 42332 27914 42334
rect 35065 42331 35131 42334
rect 16849 42256 22110 42258
rect 16849 42200 16854 42256
rect 16910 42200 22110 42256
rect 16849 42198 22110 42200
rect 16849 42195 16915 42198
rect 28206 42196 28212 42260
rect 28276 42258 28282 42260
rect 33041 42258 33107 42261
rect 28276 42256 33107 42258
rect 28276 42200 33046 42256
rect 33102 42200 33107 42256
rect 28276 42198 33107 42200
rect 28276 42196 28282 42198
rect 33041 42195 33107 42198
rect 33501 42258 33567 42261
rect 62614 42258 62620 42260
rect 33501 42256 62620 42258
rect 33501 42200 33506 42256
rect 33562 42200 62620 42256
rect 33501 42198 62620 42200
rect 33501 42195 33567 42198
rect 62614 42196 62620 42198
rect 62684 42196 62690 42260
rect 17902 42060 17908 42124
rect 17972 42122 17978 42124
rect 45553 42122 45619 42125
rect 17972 42120 45619 42122
rect 17972 42064 45558 42120
rect 45614 42064 45619 42120
rect 17972 42062 45619 42064
rect 17972 42060 17978 42062
rect 45553 42059 45619 42062
rect 27061 41986 27127 41989
rect 27705 41986 27771 41989
rect 27061 41984 27771 41986
rect 27061 41928 27066 41984
rect 27122 41928 27710 41984
rect 27766 41928 27771 41984
rect 27061 41926 27771 41928
rect 27061 41923 27127 41926
rect 27705 41923 27771 41926
rect 30373 41986 30439 41989
rect 30966 41986 30972 41988
rect 30373 41984 30972 41986
rect 30373 41928 30378 41984
rect 30434 41928 30972 41984
rect 30373 41926 30972 41928
rect 30373 41923 30439 41926
rect 30966 41924 30972 41926
rect 31036 41924 31042 41988
rect 31109 41986 31175 41989
rect 41873 41986 41939 41989
rect 31109 41984 41939 41986
rect 31109 41928 31114 41984
rect 31170 41928 41878 41984
rect 41934 41928 41939 41984
rect 31109 41926 41939 41928
rect 31109 41923 31175 41926
rect 41873 41923 41939 41926
rect 2914 41920 3230 41921
rect 2914 41856 2920 41920
rect 2984 41856 3000 41920
rect 3064 41856 3080 41920
rect 3144 41856 3160 41920
rect 3224 41856 3230 41920
rect 2914 41855 3230 41856
rect 51914 41920 52230 41921
rect 51914 41856 51920 41920
rect 51984 41856 52000 41920
rect 52064 41856 52080 41920
rect 52144 41856 52160 41920
rect 52224 41856 52230 41920
rect 51914 41855 52230 41856
rect 28717 41850 28783 41853
rect 44817 41850 44883 41853
rect 28717 41848 44883 41850
rect 28717 41792 28722 41848
rect 28778 41792 44822 41848
rect 44878 41792 44883 41848
rect 28717 41790 44883 41792
rect 28717 41787 28783 41790
rect 44817 41787 44883 41790
rect 24025 41714 24091 41717
rect 31109 41714 31175 41717
rect 36118 41714 36124 41716
rect 24025 41712 31175 41714
rect 24025 41656 24030 41712
rect 24086 41656 31114 41712
rect 31170 41656 31175 41712
rect 24025 41654 31175 41656
rect 24025 41651 24091 41654
rect 31109 41651 31175 41654
rect 31710 41654 36124 41714
rect 22369 41578 22435 41581
rect 31710 41578 31770 41654
rect 36118 41652 36124 41654
rect 36188 41652 36194 41716
rect 22369 41576 31770 41578
rect 22369 41520 22374 41576
rect 22430 41520 31770 41576
rect 22369 41518 31770 41520
rect 31845 41578 31911 41581
rect 36629 41578 36695 41581
rect 31845 41576 36695 41578
rect 31845 41520 31850 41576
rect 31906 41520 36634 41576
rect 36690 41520 36695 41576
rect 31845 41518 36695 41520
rect 22369 41515 22435 41518
rect 31845 41515 31911 41518
rect 36629 41515 36695 41518
rect 19149 41442 19215 41445
rect 27705 41442 27771 41445
rect 19149 41440 27771 41442
rect 19149 41384 19154 41440
rect 19210 41384 27710 41440
rect 27766 41384 27771 41440
rect 19149 41382 27771 41384
rect 19149 41379 19215 41382
rect 27705 41379 27771 41382
rect 34513 41442 34579 41445
rect 35014 41442 35020 41444
rect 34513 41440 35020 41442
rect 34513 41384 34518 41440
rect 34574 41384 35020 41440
rect 34513 41382 35020 41384
rect 34513 41379 34579 41382
rect 35014 41380 35020 41382
rect 35084 41380 35090 41444
rect 1994 41376 2310 41377
rect 1994 41312 2000 41376
rect 2064 41312 2080 41376
rect 2144 41312 2160 41376
rect 2224 41312 2240 41376
rect 2304 41312 2310 41376
rect 1994 41311 2310 41312
rect 50994 41376 51310 41377
rect 50994 41312 51000 41376
rect 51064 41312 51080 41376
rect 51144 41312 51160 41376
rect 51224 41312 51240 41376
rect 51304 41312 51310 41376
rect 50994 41311 51310 41312
rect 15653 41306 15719 41309
rect 26141 41306 26207 41309
rect 15653 41304 26207 41306
rect 15653 41248 15658 41304
rect 15714 41248 26146 41304
rect 26202 41248 26207 41304
rect 15653 41246 26207 41248
rect 15653 41243 15719 41246
rect 26141 41243 26207 41246
rect 26734 41244 26740 41308
rect 26804 41306 26810 41308
rect 37089 41306 37155 41309
rect 26804 41304 37155 41306
rect 26804 41248 37094 41304
rect 37150 41248 37155 41304
rect 26804 41246 37155 41248
rect 26804 41244 26810 41246
rect 37089 41243 37155 41246
rect 22134 41108 22140 41172
rect 22204 41170 22210 41172
rect 27153 41170 27219 41173
rect 34789 41170 34855 41173
rect 22204 41168 27219 41170
rect 22204 41112 27158 41168
rect 27214 41112 27219 41168
rect 22204 41110 27219 41112
rect 22204 41108 22210 41110
rect 27153 41107 27219 41110
rect 27294 41168 34855 41170
rect 27294 41112 34794 41168
rect 34850 41112 34855 41168
rect 27294 41110 34855 41112
rect 25497 41034 25563 41037
rect 27294 41034 27354 41110
rect 34789 41107 34855 41110
rect 36997 41170 37063 41173
rect 36997 41168 41430 41170
rect 36997 41112 37002 41168
rect 37058 41112 41430 41168
rect 36997 41110 41430 41112
rect 36997 41107 37063 41110
rect 25497 41032 27354 41034
rect 25497 40976 25502 41032
rect 25558 40976 27354 41032
rect 25497 40974 27354 40976
rect 25497 40971 25563 40974
rect 28942 40972 28948 41036
rect 29012 41034 29018 41036
rect 30373 41034 30439 41037
rect 29012 41032 30439 41034
rect 29012 40976 30378 41032
rect 30434 40976 30439 41032
rect 29012 40974 30439 40976
rect 29012 40972 29018 40974
rect 30373 40971 30439 40974
rect 31845 41034 31911 41037
rect 37089 41034 37155 41037
rect 31845 41032 37155 41034
rect 31845 40976 31850 41032
rect 31906 40976 37094 41032
rect 37150 40976 37155 41032
rect 31845 40974 37155 40976
rect 41370 41034 41430 41110
rect 62849 41034 62915 41037
rect 41370 41032 62915 41034
rect 41370 40976 62854 41032
rect 62910 40976 62915 41032
rect 41370 40974 62915 40976
rect 31845 40971 31911 40974
rect 37089 40971 37155 40974
rect 62849 40971 62915 40974
rect 20897 40898 20963 40901
rect 32990 40898 32996 40900
rect 20897 40896 32996 40898
rect 20897 40840 20902 40896
rect 20958 40840 32996 40896
rect 20897 40838 32996 40840
rect 20897 40835 20963 40838
rect 32990 40836 32996 40838
rect 33060 40836 33066 40900
rect 36445 40898 36511 40901
rect 50613 40898 50679 40901
rect 36445 40896 50679 40898
rect 36445 40840 36450 40896
rect 36506 40840 50618 40896
rect 50674 40840 50679 40896
rect 36445 40838 50679 40840
rect 36445 40835 36511 40838
rect 50613 40835 50679 40838
rect 2914 40832 3230 40833
rect 2914 40768 2920 40832
rect 2984 40768 3000 40832
rect 3064 40768 3080 40832
rect 3144 40768 3160 40832
rect 3224 40768 3230 40832
rect 2914 40767 3230 40768
rect 51914 40832 52230 40833
rect 51914 40768 51920 40832
rect 51984 40768 52000 40832
rect 52064 40768 52080 40832
rect 52144 40768 52160 40832
rect 52224 40768 52230 40832
rect 51914 40767 52230 40768
rect 25957 40762 26023 40765
rect 49049 40762 49115 40765
rect 25957 40760 49115 40762
rect 25957 40704 25962 40760
rect 26018 40704 49054 40760
rect 49110 40704 49115 40760
rect 25957 40702 49115 40704
rect 25957 40699 26023 40702
rect 49049 40699 49115 40702
rect 11421 40626 11487 40629
rect 24853 40626 24919 40629
rect 11421 40624 24919 40626
rect 11421 40568 11426 40624
rect 11482 40568 24858 40624
rect 24914 40568 24919 40624
rect 11421 40566 24919 40568
rect 11421 40563 11487 40566
rect 24853 40563 24919 40566
rect 27061 40626 27127 40629
rect 31661 40626 31727 40629
rect 57053 40626 57119 40629
rect 27061 40624 57119 40626
rect 27061 40568 27066 40624
rect 27122 40568 31666 40624
rect 31722 40568 57058 40624
rect 57114 40568 57119 40624
rect 27061 40566 57119 40568
rect 27061 40563 27127 40566
rect 31661 40563 31727 40566
rect 57053 40563 57119 40566
rect 29269 40490 29335 40493
rect 31201 40490 31267 40493
rect 29269 40488 31267 40490
rect 29269 40432 29274 40488
rect 29330 40432 31206 40488
rect 31262 40432 31267 40488
rect 29269 40430 31267 40432
rect 29269 40427 29335 40430
rect 31201 40427 31267 40430
rect 27705 40354 27771 40357
rect 37273 40354 37339 40357
rect 27705 40352 37339 40354
rect 27705 40296 27710 40352
rect 27766 40296 37278 40352
rect 37334 40296 37339 40352
rect 27705 40294 37339 40296
rect 27705 40291 27771 40294
rect 37273 40291 37339 40294
rect 1994 40288 2310 40289
rect 1994 40224 2000 40288
rect 2064 40224 2080 40288
rect 2144 40224 2160 40288
rect 2224 40224 2240 40288
rect 2304 40224 2310 40288
rect 1994 40223 2310 40224
rect 50994 40288 51310 40289
rect 50994 40224 51000 40288
rect 51064 40224 51080 40288
rect 51144 40224 51160 40288
rect 51224 40224 51240 40288
rect 51304 40224 51310 40288
rect 50994 40223 51310 40224
rect 29729 40218 29795 40221
rect 35801 40218 35867 40221
rect 44582 40218 44588 40220
rect 29729 40216 32322 40218
rect 29729 40160 29734 40216
rect 29790 40160 32322 40216
rect 29729 40158 32322 40160
rect 29729 40155 29795 40158
rect 32029 40084 32095 40085
rect 32029 40080 32076 40084
rect 32140 40082 32146 40084
rect 32262 40082 32322 40158
rect 35801 40216 44588 40218
rect 35801 40160 35806 40216
rect 35862 40160 44588 40216
rect 35801 40158 44588 40160
rect 35801 40155 35867 40158
rect 44582 40156 44588 40158
rect 44652 40156 44658 40220
rect 60733 40218 60799 40221
rect 63534 40218 63540 40220
rect 60733 40216 63540 40218
rect 60733 40160 60738 40216
rect 60794 40160 63540 40216
rect 60733 40158 63540 40160
rect 60733 40155 60799 40158
rect 63534 40156 63540 40158
rect 63604 40156 63610 40220
rect 37365 40082 37431 40085
rect 32029 40024 32034 40080
rect 32029 40020 32076 40024
rect 32140 40022 32186 40082
rect 32262 40080 37431 40082
rect 32262 40024 37370 40080
rect 37426 40024 37431 40080
rect 32262 40022 37431 40024
rect 32140 40020 32146 40022
rect 32029 40019 32095 40020
rect 37365 40019 37431 40022
rect 12709 39946 12775 39949
rect 57697 39946 57763 39949
rect 12709 39944 57763 39946
rect 12709 39888 12714 39944
rect 12770 39888 57702 39944
rect 57758 39888 57763 39944
rect 12709 39886 57763 39888
rect 12709 39883 12775 39886
rect 57697 39883 57763 39886
rect 19006 39748 19012 39812
rect 19076 39810 19082 39812
rect 19076 39750 31770 39810
rect 19076 39748 19082 39750
rect 2914 39744 3230 39745
rect 2914 39680 2920 39744
rect 2984 39680 3000 39744
rect 3064 39680 3080 39744
rect 3144 39680 3160 39744
rect 3224 39680 3230 39744
rect 2914 39679 3230 39680
rect 11605 39674 11671 39677
rect 28809 39674 28875 39677
rect 31710 39674 31770 39750
rect 31886 39748 31892 39812
rect 31956 39810 31962 39812
rect 32857 39810 32923 39813
rect 31956 39808 32923 39810
rect 31956 39752 32862 39808
rect 32918 39752 32923 39808
rect 31956 39750 32923 39752
rect 31956 39748 31962 39750
rect 32857 39747 32923 39750
rect 38653 39810 38719 39813
rect 46974 39810 46980 39812
rect 38653 39808 46980 39810
rect 38653 39752 38658 39808
rect 38714 39752 46980 39808
rect 38653 39750 46980 39752
rect 38653 39747 38719 39750
rect 46974 39748 46980 39750
rect 47044 39748 47050 39812
rect 51914 39744 52230 39745
rect 51914 39680 51920 39744
rect 51984 39680 52000 39744
rect 52064 39680 52080 39744
rect 52144 39680 52160 39744
rect 52224 39680 52230 39744
rect 51914 39679 52230 39680
rect 45185 39674 45251 39677
rect 45461 39674 45527 39677
rect 11605 39672 28875 39674
rect 11605 39616 11610 39672
rect 11666 39616 28814 39672
rect 28870 39616 28875 39672
rect 11605 39614 28875 39616
rect 11605 39611 11671 39614
rect 28809 39611 28875 39614
rect 28950 39614 31586 39674
rect 31710 39672 45527 39674
rect 31710 39616 45190 39672
rect 45246 39616 45466 39672
rect 45522 39616 45527 39672
rect 31710 39614 45527 39616
rect 25998 39476 26004 39540
rect 26068 39538 26074 39540
rect 28950 39538 29010 39614
rect 26068 39478 29010 39538
rect 29085 39538 29151 39541
rect 29637 39538 29703 39541
rect 29085 39536 29703 39538
rect 29085 39480 29090 39536
rect 29146 39480 29642 39536
rect 29698 39480 29703 39536
rect 29085 39478 29703 39480
rect 26068 39476 26074 39478
rect 29085 39475 29151 39478
rect 29637 39475 29703 39478
rect 30833 39538 30899 39541
rect 31334 39538 31340 39540
rect 30833 39536 31340 39538
rect 30833 39480 30838 39536
rect 30894 39480 31340 39536
rect 30833 39478 31340 39480
rect 30833 39475 30899 39478
rect 31334 39476 31340 39478
rect 31404 39476 31410 39540
rect 31526 39538 31586 39614
rect 45185 39611 45251 39614
rect 45461 39611 45527 39614
rect 49141 39674 49207 39677
rect 50521 39674 50587 39677
rect 49141 39672 50587 39674
rect 49141 39616 49146 39672
rect 49202 39616 50526 39672
rect 50582 39616 50587 39672
rect 49141 39614 50587 39616
rect 49141 39611 49207 39614
rect 50521 39611 50587 39614
rect 35249 39538 35315 39541
rect 31526 39536 35315 39538
rect 31526 39480 35254 39536
rect 35310 39480 35315 39536
rect 31526 39478 35315 39480
rect 35249 39475 35315 39478
rect 15510 39340 15516 39404
rect 15580 39402 15586 39404
rect 25957 39402 26023 39405
rect 15580 39400 26023 39402
rect 15580 39344 25962 39400
rect 26018 39344 26023 39400
rect 15580 39342 26023 39344
rect 15580 39340 15586 39342
rect 25957 39339 26023 39342
rect 28942 39340 28948 39404
rect 29012 39402 29018 39404
rect 32949 39402 33015 39405
rect 29012 39400 33015 39402
rect 29012 39344 32954 39400
rect 33010 39344 33015 39400
rect 29012 39342 33015 39344
rect 29012 39340 29018 39342
rect 32949 39339 33015 39342
rect 22502 39204 22508 39268
rect 22572 39266 22578 39268
rect 32489 39266 32555 39269
rect 22572 39264 32555 39266
rect 22572 39208 32494 39264
rect 32550 39208 32555 39264
rect 22572 39206 32555 39208
rect 22572 39204 22578 39206
rect 32489 39203 32555 39206
rect 32673 39266 32739 39269
rect 38653 39266 38719 39269
rect 32673 39264 38719 39266
rect 32673 39208 32678 39264
rect 32734 39208 38658 39264
rect 38714 39208 38719 39264
rect 32673 39206 38719 39208
rect 32673 39203 32739 39206
rect 38653 39203 38719 39206
rect 1994 39200 2310 39201
rect 1994 39136 2000 39200
rect 2064 39136 2080 39200
rect 2144 39136 2160 39200
rect 2224 39136 2240 39200
rect 2304 39136 2310 39200
rect 1994 39135 2310 39136
rect 50994 39200 51310 39201
rect 50994 39136 51000 39200
rect 51064 39136 51080 39200
rect 51144 39136 51160 39200
rect 51224 39136 51240 39200
rect 51304 39136 51310 39200
rect 50994 39135 51310 39136
rect 27286 39068 27292 39132
rect 27356 39130 27362 39132
rect 32765 39130 32831 39133
rect 27356 39128 32831 39130
rect 27356 39072 32770 39128
rect 32826 39072 32831 39128
rect 27356 39070 32831 39072
rect 27356 39068 27362 39070
rect 32765 39067 32831 39070
rect 52821 38994 52887 38997
rect 22050 38992 52887 38994
rect 22050 38936 52826 38992
rect 52882 38936 52887 38992
rect 22050 38934 52887 38936
rect 19517 38722 19583 38725
rect 22050 38722 22110 38934
rect 52821 38931 52887 38934
rect 24526 38796 24532 38860
rect 24596 38858 24602 38860
rect 27470 38858 27476 38860
rect 24596 38798 27476 38858
rect 24596 38796 24602 38798
rect 27470 38796 27476 38798
rect 27540 38796 27546 38860
rect 27797 38858 27863 38861
rect 29453 38858 29519 38861
rect 27797 38856 29519 38858
rect 27797 38800 27802 38856
rect 27858 38800 29458 38856
rect 29514 38800 29519 38856
rect 27797 38798 29519 38800
rect 27797 38795 27863 38798
rect 29453 38795 29519 38798
rect 32489 38858 32555 38861
rect 40769 38858 40835 38861
rect 32489 38856 40835 38858
rect 32489 38800 32494 38856
rect 32550 38800 40774 38856
rect 40830 38800 40835 38856
rect 32489 38798 40835 38800
rect 32489 38795 32555 38798
rect 40769 38795 40835 38798
rect 41689 38858 41755 38861
rect 43621 38858 43687 38861
rect 41689 38856 43687 38858
rect 41689 38800 41694 38856
rect 41750 38800 43626 38856
rect 43682 38800 43687 38856
rect 41689 38798 43687 38800
rect 41689 38795 41755 38798
rect 43621 38795 43687 38798
rect 44541 38858 44607 38861
rect 46657 38858 46723 38861
rect 47485 38858 47551 38861
rect 44541 38856 47551 38858
rect 44541 38800 44546 38856
rect 44602 38800 46662 38856
rect 46718 38800 47490 38856
rect 47546 38800 47551 38856
rect 44541 38798 47551 38800
rect 44541 38795 44607 38798
rect 46657 38795 46723 38798
rect 47485 38795 47551 38798
rect 19517 38720 22110 38722
rect 19517 38664 19522 38720
rect 19578 38664 22110 38720
rect 19517 38662 22110 38664
rect 24117 38722 24183 38725
rect 25681 38722 25747 38725
rect 24117 38720 25747 38722
rect 24117 38664 24122 38720
rect 24178 38664 25686 38720
rect 25742 38664 25747 38720
rect 24117 38662 25747 38664
rect 19517 38659 19583 38662
rect 24117 38659 24183 38662
rect 25681 38659 25747 38662
rect 28390 38660 28396 38724
rect 28460 38722 28466 38724
rect 31201 38722 31267 38725
rect 28460 38720 31267 38722
rect 28460 38664 31206 38720
rect 31262 38664 31267 38720
rect 28460 38662 31267 38664
rect 28460 38660 28466 38662
rect 31201 38659 31267 38662
rect 2914 38656 3230 38657
rect 2914 38592 2920 38656
rect 2984 38592 3000 38656
rect 3064 38592 3080 38656
rect 3144 38592 3160 38656
rect 3224 38592 3230 38656
rect 2914 38591 3230 38592
rect 51914 38656 52230 38657
rect 51914 38592 51920 38656
rect 51984 38592 52000 38656
rect 52064 38592 52080 38656
rect 52144 38592 52160 38656
rect 52224 38592 52230 38656
rect 51914 38591 52230 38592
rect 25129 38586 25195 38589
rect 26141 38586 26207 38589
rect 35382 38586 35388 38588
rect 25129 38584 35388 38586
rect 25129 38528 25134 38584
rect 25190 38528 26146 38584
rect 26202 38528 35388 38584
rect 25129 38526 35388 38528
rect 25129 38523 25195 38526
rect 26141 38523 26207 38526
rect 35382 38524 35388 38526
rect 35452 38524 35458 38588
rect 12065 38450 12131 38453
rect 27613 38450 27679 38453
rect 12065 38448 27679 38450
rect 12065 38392 12070 38448
rect 12126 38392 27618 38448
rect 27674 38392 27679 38448
rect 12065 38390 27679 38392
rect 12065 38387 12131 38390
rect 27613 38387 27679 38390
rect 21398 38252 21404 38316
rect 21468 38314 21474 38316
rect 29545 38314 29611 38317
rect 21468 38312 29611 38314
rect 21468 38256 29550 38312
rect 29606 38256 29611 38312
rect 21468 38254 29611 38256
rect 21468 38252 21474 38254
rect 29545 38251 29611 38254
rect 32990 38252 32996 38316
rect 33060 38314 33066 38316
rect 34145 38314 34211 38317
rect 33060 38312 34211 38314
rect 33060 38256 34150 38312
rect 34206 38256 34211 38312
rect 33060 38254 34211 38256
rect 33060 38252 33066 38254
rect 34145 38251 34211 38254
rect 34421 38314 34487 38317
rect 63217 38314 63283 38317
rect 34421 38312 63283 38314
rect 34421 38256 34426 38312
rect 34482 38256 63222 38312
rect 63278 38256 63283 38312
rect 34421 38254 63283 38256
rect 34421 38251 34487 38254
rect 63217 38251 63283 38254
rect 34329 38178 34395 38181
rect 22050 38176 34395 38178
rect 22050 38120 34334 38176
rect 34390 38120 34395 38176
rect 22050 38118 34395 38120
rect 1994 38112 2310 38113
rect 1994 38048 2000 38112
rect 2064 38048 2080 38112
rect 2144 38048 2160 38112
rect 2224 38048 2240 38112
rect 2304 38048 2310 38112
rect 1994 38047 2310 38048
rect 14406 37980 14412 38044
rect 14476 38042 14482 38044
rect 22050 38042 22110 38118
rect 34329 38115 34395 38118
rect 50994 38112 51310 38113
rect 50994 38048 51000 38112
rect 51064 38048 51080 38112
rect 51144 38048 51160 38112
rect 51224 38048 51240 38112
rect 51304 38048 51310 38112
rect 50994 38047 51310 38048
rect 14476 37982 22110 38042
rect 14476 37980 14482 37982
rect 24894 37980 24900 38044
rect 24964 38042 24970 38044
rect 38009 38042 38075 38045
rect 38929 38042 38995 38045
rect 24964 38040 38995 38042
rect 24964 37984 38014 38040
rect 38070 37984 38934 38040
rect 38990 37984 38995 38040
rect 24964 37982 38995 37984
rect 24964 37980 24970 37982
rect 38009 37979 38075 37982
rect 38929 37979 38995 37982
rect 27470 37844 27476 37908
rect 27540 37906 27546 37908
rect 30230 37906 30236 37908
rect 27540 37846 30236 37906
rect 27540 37844 27546 37846
rect 30230 37844 30236 37846
rect 30300 37844 30306 37908
rect 32070 37844 32076 37908
rect 32140 37906 32146 37908
rect 32990 37906 32996 37908
rect 32140 37846 32996 37906
rect 32140 37844 32146 37846
rect 32990 37844 32996 37846
rect 33060 37844 33066 37908
rect 33133 37906 33199 37909
rect 50061 37906 50127 37909
rect 33133 37904 50127 37906
rect 33133 37848 33138 37904
rect 33194 37848 50066 37904
rect 50122 37848 50127 37904
rect 33133 37846 50127 37848
rect 33133 37843 33199 37846
rect 50061 37843 50127 37846
rect 14825 37770 14891 37773
rect 55397 37770 55463 37773
rect 55857 37770 55923 37773
rect 14825 37768 55923 37770
rect 14825 37712 14830 37768
rect 14886 37712 55402 37768
rect 55458 37712 55862 37768
rect 55918 37712 55923 37768
rect 14825 37710 55923 37712
rect 14825 37707 14891 37710
rect 55397 37707 55463 37710
rect 55857 37707 55923 37710
rect 20110 37572 20116 37636
rect 20180 37634 20186 37636
rect 43805 37634 43871 37637
rect 20180 37632 43871 37634
rect 20180 37576 43810 37632
rect 43866 37576 43871 37632
rect 20180 37574 43871 37576
rect 20180 37572 20186 37574
rect 43805 37571 43871 37574
rect 2914 37568 3230 37569
rect 2914 37504 2920 37568
rect 2984 37504 3000 37568
rect 3064 37504 3080 37568
rect 3144 37504 3160 37568
rect 3224 37504 3230 37568
rect 2914 37503 3230 37504
rect 51914 37568 52230 37569
rect 51914 37504 51920 37568
rect 51984 37504 52000 37568
rect 52064 37504 52080 37568
rect 52144 37504 52160 37568
rect 52224 37504 52230 37568
rect 51914 37503 52230 37504
rect 65254 37568 65570 37569
rect 65254 37504 65260 37568
rect 65324 37504 65340 37568
rect 65404 37504 65420 37568
rect 65484 37504 65500 37568
rect 65564 37504 65570 37568
rect 65254 37503 65570 37504
rect 29310 37436 29316 37500
rect 29380 37498 29386 37500
rect 34513 37498 34579 37501
rect 29380 37496 34579 37498
rect 29380 37440 34518 37496
rect 34574 37440 34579 37496
rect 29380 37438 34579 37440
rect 29380 37436 29386 37438
rect 34513 37435 34579 37438
rect 15101 37362 15167 37365
rect 27889 37362 27955 37365
rect 15101 37360 27955 37362
rect 15101 37304 15106 37360
rect 15162 37304 27894 37360
rect 27950 37304 27955 37360
rect 15101 37302 27955 37304
rect 15101 37299 15167 37302
rect 27889 37299 27955 37302
rect 28533 37362 28599 37365
rect 33685 37364 33751 37365
rect 32070 37362 32076 37364
rect 28533 37360 32076 37362
rect 28533 37304 28538 37360
rect 28594 37304 32076 37360
rect 28533 37302 32076 37304
rect 28533 37299 28599 37302
rect 32070 37300 32076 37302
rect 32140 37300 32146 37364
rect 32262 37302 32690 37362
rect 21633 37226 21699 37229
rect 32262 37226 32322 37302
rect 21633 37224 32322 37226
rect 21633 37168 21638 37224
rect 21694 37168 32322 37224
rect 21633 37166 32322 37168
rect 32397 37228 32463 37229
rect 32397 37224 32444 37228
rect 32508 37226 32514 37228
rect 32630 37226 32690 37302
rect 33685 37360 33732 37364
rect 33796 37362 33802 37364
rect 35801 37362 35867 37365
rect 62021 37362 62087 37365
rect 33685 37304 33690 37360
rect 33685 37300 33732 37304
rect 33796 37302 33842 37362
rect 35801 37360 62087 37362
rect 35801 37304 35806 37360
rect 35862 37304 62026 37360
rect 62082 37304 62087 37360
rect 35801 37302 62087 37304
rect 33796 37300 33802 37302
rect 33685 37299 33751 37300
rect 35801 37299 35867 37302
rect 62021 37299 62087 37302
rect 33358 37226 33364 37228
rect 32397 37168 32402 37224
rect 21633 37163 21699 37166
rect 32397 37164 32444 37168
rect 32508 37166 32554 37226
rect 32630 37166 33364 37226
rect 32508 37164 32514 37166
rect 33358 37164 33364 37166
rect 33428 37164 33434 37228
rect 34421 37226 34487 37229
rect 42374 37226 42380 37228
rect 34421 37224 42380 37226
rect 34421 37168 34426 37224
rect 34482 37168 42380 37224
rect 34421 37166 42380 37168
rect 32397 37163 32463 37164
rect 34421 37163 34487 37166
rect 42374 37164 42380 37166
rect 42444 37164 42450 37228
rect 10910 37028 10916 37092
rect 10980 37090 10986 37092
rect 19517 37090 19583 37093
rect 10980 37088 19583 37090
rect 10980 37032 19522 37088
rect 19578 37032 19583 37088
rect 10980 37030 19583 37032
rect 10980 37028 10986 37030
rect 19517 37027 19583 37030
rect 21030 37028 21036 37092
rect 21100 37090 21106 37092
rect 26049 37090 26115 37093
rect 21100 37088 26115 37090
rect 21100 37032 26054 37088
rect 26110 37032 26115 37088
rect 21100 37030 26115 37032
rect 21100 37028 21106 37030
rect 26049 37027 26115 37030
rect 29085 37090 29151 37093
rect 32806 37090 32812 37092
rect 29085 37088 32812 37090
rect 29085 37032 29090 37088
rect 29146 37032 32812 37088
rect 29085 37030 32812 37032
rect 29085 37027 29151 37030
rect 32806 37028 32812 37030
rect 32876 37028 32882 37092
rect 1994 37024 2310 37025
rect 1994 36960 2000 37024
rect 2064 36960 2080 37024
rect 2144 36960 2160 37024
rect 2224 36960 2240 37024
rect 2304 36960 2310 37024
rect 1994 36959 2310 36960
rect 50994 37024 51310 37025
rect 50994 36960 51000 37024
rect 51064 36960 51080 37024
rect 51144 36960 51160 37024
rect 51224 36960 51240 37024
rect 51304 36960 51310 37024
rect 50994 36959 51310 36960
rect 64334 37024 64650 37025
rect 64334 36960 64340 37024
rect 64404 36960 64420 37024
rect 64484 36960 64500 37024
rect 64564 36960 64580 37024
rect 64644 36960 64650 37024
rect 64334 36959 64650 36960
rect 9622 36892 9628 36956
rect 9692 36954 9698 36956
rect 20345 36954 20411 36957
rect 21633 36956 21699 36957
rect 21582 36954 21588 36956
rect 9692 36952 20411 36954
rect 9692 36896 20350 36952
rect 20406 36896 20411 36952
rect 9692 36894 20411 36896
rect 21542 36894 21588 36954
rect 21652 36952 21699 36956
rect 21694 36896 21699 36952
rect 9692 36892 9698 36894
rect 20345 36891 20411 36894
rect 21582 36892 21588 36894
rect 21652 36892 21699 36896
rect 23790 36892 23796 36956
rect 23860 36954 23866 36956
rect 36813 36954 36879 36957
rect 23860 36952 36879 36954
rect 23860 36896 36818 36952
rect 36874 36896 36879 36952
rect 23860 36894 36879 36896
rect 23860 36892 23866 36894
rect 21633 36891 21699 36892
rect 36813 36891 36879 36894
rect 12014 36756 12020 36820
rect 12084 36818 12090 36820
rect 23197 36818 23263 36821
rect 12084 36816 23263 36818
rect 12084 36760 23202 36816
rect 23258 36760 23263 36816
rect 12084 36758 23263 36760
rect 12084 36756 12090 36758
rect 23197 36755 23263 36758
rect 24761 36818 24827 36821
rect 30373 36818 30439 36821
rect 24761 36816 30439 36818
rect 24761 36760 24766 36816
rect 24822 36760 30378 36816
rect 30434 36760 30439 36816
rect 24761 36758 30439 36760
rect 24761 36755 24827 36758
rect 30373 36755 30439 36758
rect 30598 36756 30604 36820
rect 30668 36818 30674 36820
rect 45870 36818 45876 36820
rect 30668 36758 45876 36818
rect 30668 36756 30674 36758
rect 45870 36756 45876 36758
rect 45940 36756 45946 36820
rect 6126 36620 6132 36684
rect 6196 36682 6202 36684
rect 15101 36682 15167 36685
rect 6196 36680 15167 36682
rect 6196 36624 15106 36680
rect 15162 36624 15167 36680
rect 6196 36622 15167 36624
rect 6196 36620 6202 36622
rect 15101 36619 15167 36622
rect 15285 36682 15351 36685
rect 39982 36682 39988 36684
rect 15285 36680 39988 36682
rect 15285 36624 15290 36680
rect 15346 36624 39988 36680
rect 15285 36622 39988 36624
rect 15285 36619 15351 36622
rect 39982 36620 39988 36622
rect 40052 36620 40058 36684
rect 66529 36682 66595 36685
rect 41370 36680 66595 36682
rect 41370 36624 66534 36680
rect 66590 36624 66595 36680
rect 41370 36622 66595 36624
rect 3918 36484 3924 36548
rect 3988 36546 3994 36548
rect 23606 36546 23612 36548
rect 3988 36486 23612 36546
rect 3988 36484 3994 36486
rect 23606 36484 23612 36486
rect 23676 36484 23682 36548
rect 30097 36546 30163 36549
rect 41370 36546 41430 36622
rect 66529 36619 66595 36622
rect 30097 36544 41430 36546
rect 30097 36488 30102 36544
rect 30158 36488 41430 36544
rect 30097 36486 41430 36488
rect 30097 36483 30163 36486
rect 65254 36480 65570 36481
rect 65254 36416 65260 36480
rect 65324 36416 65340 36480
rect 65404 36416 65420 36480
rect 65484 36416 65500 36480
rect 65564 36416 65570 36480
rect 65254 36415 65570 36416
rect 25078 36348 25084 36412
rect 25148 36410 25154 36412
rect 30465 36410 30531 36413
rect 25148 36408 30531 36410
rect 25148 36352 30470 36408
rect 30526 36352 30531 36408
rect 25148 36350 30531 36352
rect 25148 36348 25154 36350
rect 30465 36347 30531 36350
rect 32857 36410 32923 36413
rect 64086 36410 64092 36412
rect 32857 36408 64092 36410
rect 32857 36352 32862 36408
rect 32918 36352 64092 36408
rect 32857 36350 64092 36352
rect 32857 36347 32923 36350
rect 64086 36348 64092 36350
rect 64156 36348 64162 36412
rect 19558 36212 19564 36276
rect 19628 36274 19634 36276
rect 24025 36274 24091 36277
rect 19628 36272 24091 36274
rect 19628 36216 24030 36272
rect 24086 36216 24091 36272
rect 19628 36214 24091 36216
rect 19628 36212 19634 36214
rect 24025 36211 24091 36214
rect 28993 36274 29059 36277
rect 37273 36274 37339 36277
rect 62573 36274 62639 36277
rect 28993 36272 34346 36274
rect 28993 36216 28998 36272
rect 29054 36216 34346 36272
rect 28993 36214 34346 36216
rect 28993 36211 29059 36214
rect 16614 36076 16620 36140
rect 16684 36138 16690 36140
rect 25497 36138 25563 36141
rect 16684 36136 25563 36138
rect 16684 36080 25502 36136
rect 25558 36080 25563 36136
rect 16684 36078 25563 36080
rect 16684 36076 16690 36078
rect 25497 36075 25563 36078
rect 4976 35940 4982 36004
rect 5046 36002 5052 36004
rect 12157 36002 12223 36005
rect 5046 36000 12223 36002
rect 5046 35944 12162 36000
rect 12218 35944 12223 36000
rect 5046 35942 12223 35944
rect 5046 35940 5052 35942
rect 12157 35939 12223 35942
rect 13152 35940 13158 36004
rect 13222 36002 13228 36004
rect 19701 36002 19767 36005
rect 13222 36000 19767 36002
rect 13222 35944 19706 36000
rect 19762 35944 19767 36000
rect 13222 35942 19767 35944
rect 13222 35940 13228 35942
rect 19701 35939 19767 35942
rect 26468 35940 26474 36004
rect 26538 36002 26544 36004
rect 31661 36002 31727 36005
rect 26538 36000 31727 36002
rect 26538 35944 31666 36000
rect 31722 35944 31727 36000
rect 26538 35942 31727 35944
rect 26538 35940 26544 35942
rect 31661 35939 31727 35942
rect 33409 36002 33475 36005
rect 34038 36002 34044 36004
rect 33409 36000 34044 36002
rect 33409 35944 33414 36000
rect 33470 35944 34044 36000
rect 33409 35942 34044 35944
rect 33409 35939 33475 35942
rect 34038 35940 34044 35942
rect 34108 35940 34114 36004
rect 34286 36002 34346 36214
rect 37273 36272 62639 36274
rect 37273 36216 37278 36272
rect 37334 36216 62578 36272
rect 62634 36216 62639 36272
rect 37273 36214 62639 36216
rect 37273 36211 37339 36214
rect 62573 36211 62639 36214
rect 63585 36274 63651 36277
rect 63902 36274 63908 36276
rect 63585 36272 63908 36274
rect 63585 36216 63590 36272
rect 63646 36216 63908 36272
rect 63585 36214 63908 36216
rect 63585 36211 63651 36214
rect 63902 36212 63908 36214
rect 63972 36212 63978 36276
rect 34421 36138 34487 36141
rect 62665 36138 62731 36141
rect 34421 36136 62731 36138
rect 34421 36080 34426 36136
rect 34482 36080 62670 36136
rect 62726 36080 62731 36136
rect 34421 36078 62731 36080
rect 34421 36075 34487 36078
rect 62665 36075 62731 36078
rect 37680 36002 37686 36004
rect 34286 35942 37686 36002
rect 37680 35940 37686 35942
rect 37750 35940 37756 36004
rect 62113 36002 62179 36005
rect 63350 36002 63356 36004
rect 62113 36000 63356 36002
rect 62113 35944 62118 36000
rect 62174 35944 63356 36000
rect 62113 35942 63356 35944
rect 62113 35939 62179 35942
rect 63350 35940 63356 35942
rect 63420 35940 63426 36004
rect 64334 35936 64650 35937
rect 64334 35872 64340 35936
rect 64404 35872 64420 35936
rect 64484 35872 64500 35936
rect 64564 35872 64580 35936
rect 64644 35872 64650 35936
rect 64334 35871 64650 35872
rect 22001 35868 22067 35869
rect 23565 35868 23631 35869
rect 24485 35868 24551 35869
rect 24761 35868 24827 35869
rect 25865 35868 25931 35869
rect 21962 35866 21968 35868
rect 21910 35806 21968 35866
rect 22032 35864 22067 35868
rect 23526 35866 23532 35868
rect 22062 35808 22067 35864
rect 21962 35804 21968 35806
rect 22032 35804 22067 35808
rect 23474 35806 23532 35866
rect 23596 35864 23631 35868
rect 24468 35866 24474 35868
rect 23626 35808 23631 35864
rect 23526 35804 23532 35806
rect 23596 35804 23631 35808
rect 24394 35806 24474 35866
rect 24538 35864 24551 35868
rect 24546 35808 24551 35864
rect 24468 35804 24474 35806
rect 24538 35804 24551 35808
rect 24710 35804 24716 35868
rect 24780 35866 24827 35868
rect 24780 35864 24872 35866
rect 24822 35808 24872 35864
rect 24780 35806 24872 35808
rect 24780 35804 24827 35806
rect 25862 35804 25868 35868
rect 25932 35866 25938 35868
rect 25932 35806 26022 35866
rect 25932 35804 25938 35806
rect 29504 35804 29510 35868
rect 29574 35866 29580 35868
rect 30005 35866 30071 35869
rect 29574 35864 30071 35866
rect 29574 35808 30010 35864
rect 30066 35808 30071 35864
rect 29574 35806 30071 35808
rect 29574 35804 29580 35806
rect 22001 35803 22067 35804
rect 23565 35803 23631 35804
rect 24485 35803 24551 35804
rect 24761 35803 24827 35804
rect 25865 35803 25931 35804
rect 30005 35803 30071 35806
rect 30189 35868 30255 35869
rect 30189 35864 30198 35868
rect 30262 35866 30268 35868
rect 30189 35808 30194 35864
rect 30189 35804 30198 35808
rect 30262 35806 30346 35866
rect 30262 35804 30268 35806
rect 30690 35804 30696 35868
rect 30760 35866 30766 35868
rect 31109 35866 31175 35869
rect 31840 35866 31846 35868
rect 30760 35864 31175 35866
rect 30760 35808 31114 35864
rect 31170 35808 31175 35864
rect 30760 35806 31175 35808
rect 30760 35804 30766 35806
rect 30189 35803 30255 35804
rect 31109 35803 31175 35806
rect 31710 35806 31846 35866
rect 7322 35668 7328 35732
rect 7392 35730 7398 35732
rect 8201 35730 8267 35733
rect 7392 35728 8267 35730
rect 7392 35672 8206 35728
rect 8262 35672 8267 35728
rect 7392 35670 8267 35672
rect 7392 35668 7398 35670
rect 8201 35667 8267 35670
rect 8480 35668 8486 35732
rect 8550 35730 8556 35732
rect 15009 35730 15075 35733
rect 20069 35732 20135 35733
rect 20022 35730 20028 35732
rect 8550 35728 15075 35730
rect 8550 35672 15014 35728
rect 15070 35672 15075 35728
rect 8550 35670 15075 35672
rect 19978 35670 20028 35730
rect 20092 35728 20135 35732
rect 20130 35672 20135 35728
rect 8550 35668 8556 35670
rect 15009 35667 15075 35670
rect 20022 35668 20028 35670
rect 20092 35668 20135 35672
rect 21190 35668 21196 35732
rect 21260 35730 21266 35732
rect 21357 35730 21423 35733
rect 21260 35728 21423 35730
rect 21260 35672 21362 35728
rect 21418 35672 21423 35728
rect 21260 35670 21423 35672
rect 21260 35668 21266 35670
rect 20069 35667 20135 35668
rect 21357 35667 21423 35670
rect 22185 35732 22251 35733
rect 23013 35732 23079 35733
rect 23197 35732 23263 35733
rect 25221 35732 25287 35733
rect 22185 35728 22198 35732
rect 22262 35730 22268 35732
rect 22962 35730 22968 35732
rect 22185 35672 22190 35728
rect 22185 35668 22198 35672
rect 22262 35670 22342 35730
rect 22922 35670 22968 35730
rect 23032 35728 23079 35732
rect 23074 35672 23079 35728
rect 22262 35668 22268 35670
rect 22962 35668 22968 35670
rect 23032 35668 23079 35672
rect 23192 35668 23198 35732
rect 23262 35730 23268 35732
rect 25204 35730 25210 35732
rect 23262 35670 23350 35730
rect 25130 35670 25210 35730
rect 25274 35728 25287 35732
rect 25282 35672 25287 35728
rect 23262 35668 23268 35670
rect 25204 35668 25210 35670
rect 25274 35668 25287 35672
rect 29962 35668 29968 35732
rect 30032 35730 30038 35732
rect 30281 35730 30347 35733
rect 30032 35728 30347 35730
rect 30032 35672 30286 35728
rect 30342 35672 30347 35728
rect 30032 35670 30347 35672
rect 30032 35668 30038 35670
rect 22185 35667 22251 35668
rect 23013 35667 23079 35668
rect 23197 35667 23263 35668
rect 25221 35667 25287 35668
rect 30281 35667 30347 35670
rect 30465 35730 30531 35733
rect 31710 35730 31770 35806
rect 31840 35804 31846 35806
rect 31910 35804 31916 35868
rect 33041 35866 33107 35869
rect 34176 35866 34182 35868
rect 33041 35864 34182 35866
rect 33041 35808 33046 35864
rect 33102 35808 34182 35864
rect 33041 35806 34182 35808
rect 33041 35803 33107 35806
rect 34176 35804 34182 35806
rect 34246 35804 34252 35868
rect 34513 35866 34579 35869
rect 35192 35866 35198 35868
rect 34513 35864 35198 35866
rect 34513 35808 34518 35864
rect 34574 35808 35198 35864
rect 34513 35806 35198 35808
rect 34513 35803 34579 35806
rect 35192 35804 35198 35806
rect 35262 35804 35268 35868
rect 38561 35866 38627 35869
rect 38848 35866 38854 35868
rect 38561 35864 38854 35866
rect 38561 35808 38566 35864
rect 38622 35808 38854 35864
rect 38561 35806 38854 35808
rect 38561 35803 38627 35806
rect 38848 35804 38854 35806
rect 38918 35804 38924 35868
rect 42701 35866 42767 35869
rect 43520 35866 43526 35868
rect 42701 35864 43526 35866
rect 42701 35808 42706 35864
rect 42762 35808 43526 35864
rect 42701 35806 43526 35808
rect 42701 35803 42767 35806
rect 43520 35804 43526 35806
rect 43590 35804 43596 35868
rect 36537 35732 36603 35733
rect 36512 35730 36518 35732
rect 30465 35728 31770 35730
rect 30465 35672 30470 35728
rect 30526 35672 31770 35728
rect 30465 35670 31770 35672
rect 36446 35670 36518 35730
rect 36582 35728 36603 35732
rect 36598 35672 36603 35728
rect 30465 35667 30531 35670
rect 36512 35668 36518 35670
rect 36582 35668 36603 35672
rect 36537 35667 36603 35668
rect 38653 35730 38719 35733
rect 41178 35730 41184 35732
rect 38653 35728 41184 35730
rect 38653 35672 38658 35728
rect 38714 35672 41184 35728
rect 38653 35670 41184 35672
rect 38653 35667 38719 35670
rect 41178 35668 41184 35670
rect 41248 35668 41254 35732
rect 56240 35668 56246 35732
rect 56310 35730 56316 35732
rect 56409 35730 56475 35733
rect 63953 35730 64019 35733
rect 56310 35728 64019 35730
rect 56310 35672 56414 35728
rect 56470 35672 63958 35728
rect 64014 35672 64019 35728
rect 56310 35670 64019 35672
rect 56310 35668 56316 35670
rect 56409 35667 56475 35670
rect 63953 35667 64019 35670
rect 1992 35492 2312 35514
rect 1992 35428 2000 35492
rect 2064 35428 2080 35492
rect 2144 35428 2160 35492
rect 2224 35428 2240 35492
rect 2304 35428 2312 35492
rect 1992 35412 2312 35428
rect 1992 35348 2000 35412
rect 2064 35348 2080 35412
rect 2144 35348 2160 35412
rect 2224 35348 2240 35412
rect 2304 35348 2312 35412
rect 1992 35332 2312 35348
rect 1992 35268 2000 35332
rect 2064 35268 2080 35332
rect 2144 35268 2160 35332
rect 2224 35268 2240 35332
rect 2304 35268 2312 35332
rect 1992 35252 2312 35268
rect 1992 35188 2000 35252
rect 2064 35188 2080 35252
rect 2144 35188 2160 35252
rect 2224 35188 2240 35252
rect 2304 35188 2312 35252
rect 1992 35166 2312 35188
rect 50992 35492 51312 35514
rect 50992 35428 51000 35492
rect 51064 35428 51080 35492
rect 51144 35428 51160 35492
rect 51224 35428 51240 35492
rect 51304 35428 51312 35492
rect 50992 35412 51312 35428
rect 50992 35348 51000 35412
rect 51064 35348 51080 35412
rect 51144 35348 51160 35412
rect 51224 35348 51240 35412
rect 51304 35348 51312 35412
rect 50992 35332 51312 35348
rect 50992 35268 51000 35332
rect 51064 35268 51080 35332
rect 51144 35268 51160 35332
rect 51224 35268 51240 35332
rect 51304 35268 51312 35332
rect 65254 35392 65570 35393
rect 65254 35328 65260 35392
rect 65324 35328 65340 35392
rect 65404 35328 65420 35392
rect 65484 35328 65500 35392
rect 65564 35328 65570 35392
rect 65254 35327 65570 35328
rect 50992 35252 51312 35268
rect 50992 35188 51000 35252
rect 51064 35188 51080 35252
rect 51144 35188 51160 35252
rect 51224 35188 51240 35252
rect 51304 35188 51312 35252
rect 50992 35166 51312 35188
rect 64334 34848 64650 34849
rect 2912 34796 3232 34818
rect 2912 34732 2920 34796
rect 2984 34732 3000 34796
rect 3064 34732 3080 34796
rect 3144 34732 3160 34796
rect 3224 34732 3232 34796
rect 2912 34716 3232 34732
rect 2912 34652 2920 34716
rect 2984 34652 3000 34716
rect 3064 34652 3080 34716
rect 3144 34652 3160 34716
rect 3224 34652 3232 34716
rect 2912 34636 3232 34652
rect 2912 34572 2920 34636
rect 2984 34572 3000 34636
rect 3064 34572 3080 34636
rect 3144 34572 3160 34636
rect 3224 34572 3232 34636
rect 2912 34556 3232 34572
rect 2912 34492 2920 34556
rect 2984 34492 3000 34556
rect 3064 34492 3080 34556
rect 3144 34492 3160 34556
rect 3224 34492 3232 34556
rect 2912 34470 3232 34492
rect 51912 34796 52232 34818
rect 51912 34732 51920 34796
rect 51984 34732 52000 34796
rect 52064 34732 52080 34796
rect 52144 34732 52160 34796
rect 52224 34732 52232 34796
rect 64334 34784 64340 34848
rect 64404 34784 64420 34848
rect 64484 34784 64500 34848
rect 64564 34784 64580 34848
rect 64644 34784 64650 34848
rect 64334 34783 64650 34784
rect 51912 34716 52232 34732
rect 51912 34652 51920 34716
rect 51984 34652 52000 34716
rect 52064 34652 52080 34716
rect 52144 34652 52160 34716
rect 52224 34652 52232 34716
rect 63493 34778 63559 34781
rect 63718 34778 63724 34780
rect 63493 34776 63724 34778
rect 63493 34720 63498 34776
rect 63554 34720 63724 34776
rect 63493 34718 63724 34720
rect 63493 34715 63559 34718
rect 63718 34716 63724 34718
rect 63788 34716 63794 34780
rect 51912 34636 52232 34652
rect 51912 34572 51920 34636
rect 51984 34572 52000 34636
rect 52064 34572 52080 34636
rect 52144 34572 52160 34636
rect 52224 34572 52232 34636
rect 63534 34580 63540 34644
rect 63604 34642 63610 34644
rect 63677 34642 63743 34645
rect 63604 34640 63743 34642
rect 63604 34584 63682 34640
rect 63738 34584 63743 34640
rect 63604 34582 63743 34584
rect 63604 34580 63610 34582
rect 63677 34579 63743 34582
rect 51912 34556 52232 34572
rect 51912 34492 51920 34556
rect 51984 34492 52000 34556
rect 52064 34492 52080 34556
rect 52144 34492 52160 34556
rect 52224 34492 52232 34556
rect 51912 34470 52232 34492
rect 65254 34304 65570 34305
rect 65254 34240 65260 34304
rect 65324 34240 65340 34304
rect 65404 34240 65420 34304
rect 65484 34240 65500 34304
rect 65564 34240 65570 34304
rect 65254 34239 65570 34240
rect 64334 33760 64650 33761
rect 64334 33696 64340 33760
rect 64404 33696 64420 33760
rect 64484 33696 64500 33760
rect 64564 33696 64580 33760
rect 64644 33696 64650 33760
rect 64334 33695 64650 33696
rect 65254 33216 65570 33217
rect 65254 33152 65260 33216
rect 65324 33152 65340 33216
rect 65404 33152 65420 33216
rect 65484 33152 65500 33216
rect 65564 33152 65570 33216
rect 65254 33151 65570 33152
rect 64334 32672 64650 32673
rect 64334 32608 64340 32672
rect 64404 32608 64420 32672
rect 64484 32608 64500 32672
rect 64564 32608 64580 32672
rect 64644 32608 64650 32672
rect 64334 32607 64650 32608
rect 65254 32128 65570 32129
rect 65254 32064 65260 32128
rect 65324 32064 65340 32128
rect 65404 32064 65420 32128
rect 65484 32064 65500 32128
rect 65564 32064 65570 32128
rect 65254 32063 65570 32064
rect 64334 31584 64650 31585
rect 64334 31520 64340 31584
rect 64404 31520 64420 31584
rect 64484 31520 64500 31584
rect 64564 31520 64580 31584
rect 64644 31520 64650 31584
rect 64334 31519 64650 31520
rect 62665 31240 62731 31245
rect 62665 31184 62670 31240
rect 62726 31184 62731 31240
rect 62665 31179 62731 31184
rect 62668 30940 62728 31179
rect 65254 31040 65570 31041
rect 65254 30976 65260 31040
rect 65324 30976 65340 31040
rect 65404 30976 65420 31040
rect 65484 30976 65500 31040
rect 65564 30976 65570 31040
rect 65254 30975 65570 30976
rect 62504 30880 62728 30940
rect 64334 30496 64650 30497
rect 64334 30432 64340 30496
rect 64404 30432 64420 30496
rect 64484 30432 64500 30496
rect 64564 30432 64580 30496
rect 64644 30432 64650 30496
rect 64334 30431 64650 30432
rect 65254 29952 65570 29953
rect 65254 29888 65260 29952
rect 65324 29888 65340 29952
rect 65404 29888 65420 29952
rect 65484 29888 65500 29952
rect 65564 29888 65570 29952
rect 65254 29887 65570 29888
rect 64334 29408 64650 29409
rect 64334 29344 64340 29408
rect 64404 29344 64420 29408
rect 64484 29344 64500 29408
rect 64564 29344 64580 29408
rect 64644 29344 64650 29408
rect 64334 29343 64650 29344
rect 62614 29240 62620 29242
rect 62504 29180 62620 29240
rect 62614 29178 62620 29180
rect 62684 29178 62690 29242
rect 64965 29066 65031 29069
rect 64830 29064 65031 29066
rect 64830 29008 64970 29064
rect 65026 29008 65031 29064
rect 64830 29006 65031 29008
rect 64830 28797 64890 29006
rect 64965 29003 65031 29006
rect 65254 28864 65570 28865
rect 65254 28800 65260 28864
rect 65324 28800 65340 28864
rect 65404 28800 65420 28864
rect 65484 28800 65500 28864
rect 65564 28800 65570 28864
rect 65254 28799 65570 28800
rect 64830 28792 64939 28797
rect 64830 28736 64878 28792
rect 64934 28736 64939 28792
rect 64830 28734 64939 28736
rect 64873 28731 64939 28734
rect 64334 28320 64650 28321
rect 64334 28256 64340 28320
rect 64404 28256 64420 28320
rect 64484 28256 64500 28320
rect 64564 28256 64580 28320
rect 64644 28256 64650 28320
rect 64334 28255 64650 28256
rect 65254 27776 65570 27777
rect 65254 27712 65260 27776
rect 65324 27712 65340 27776
rect 65404 27712 65420 27776
rect 65484 27712 65500 27776
rect 65564 27712 65570 27776
rect 65254 27711 65570 27712
rect 64334 27232 64650 27233
rect 64334 27168 64340 27232
rect 64404 27168 64420 27232
rect 64484 27168 64500 27232
rect 64564 27168 64580 27232
rect 64644 27168 64650 27232
rect 64334 27167 64650 27168
rect 65254 26688 65570 26689
rect 65254 26624 65260 26688
rect 65324 26624 65340 26688
rect 65404 26624 65420 26688
rect 65484 26624 65500 26688
rect 65564 26624 65570 26688
rect 65254 26623 65570 26624
rect 64334 26144 64650 26145
rect 64334 26080 64340 26144
rect 64404 26080 64420 26144
rect 64484 26080 64500 26144
rect 64564 26080 64580 26144
rect 64644 26080 64650 26144
rect 64334 26079 64650 26080
rect 65254 25600 65570 25601
rect 65254 25536 65260 25600
rect 65324 25536 65340 25600
rect 65404 25536 65420 25600
rect 65484 25536 65500 25600
rect 65564 25536 65570 25600
rect 65254 25535 65570 25536
rect 64334 25056 64650 25057
rect 64334 24992 64340 25056
rect 64404 24992 64420 25056
rect 64484 24992 64500 25056
rect 64564 24992 64580 25056
rect 64644 24992 64650 25056
rect 64334 24991 64650 24992
rect 65254 24512 65570 24513
rect 65254 24448 65260 24512
rect 65324 24448 65340 24512
rect 65404 24448 65420 24512
rect 65484 24448 65500 24512
rect 65564 24448 65570 24512
rect 65254 24447 65570 24448
rect 64334 23968 64650 23969
rect 64334 23904 64340 23968
rect 64404 23904 64420 23968
rect 64484 23904 64500 23968
rect 64564 23904 64580 23968
rect 64644 23904 64650 23968
rect 64334 23903 64650 23904
rect 65254 23424 65570 23425
rect 65254 23360 65260 23424
rect 65324 23360 65340 23424
rect 65404 23360 65420 23424
rect 65484 23360 65500 23424
rect 65564 23360 65570 23424
rect 65254 23359 65570 23360
rect 64334 22880 64650 22881
rect 64334 22816 64340 22880
rect 64404 22816 64420 22880
rect 64484 22816 64500 22880
rect 64564 22816 64580 22880
rect 64644 22816 64650 22880
rect 64334 22815 64650 22816
rect 65254 22336 65570 22337
rect 65254 22272 65260 22336
rect 65324 22272 65340 22336
rect 65404 22272 65420 22336
rect 65484 22272 65500 22336
rect 65564 22272 65570 22336
rect 65254 22271 65570 22272
rect 64334 21792 64650 21793
rect 64334 21728 64340 21792
rect 64404 21728 64420 21792
rect 64484 21728 64500 21792
rect 64564 21728 64580 21792
rect 64644 21728 64650 21792
rect 64334 21727 64650 21728
rect 65254 21248 65570 21249
rect 65254 21184 65260 21248
rect 65324 21184 65340 21248
rect 65404 21184 65420 21248
rect 65484 21184 65500 21248
rect 65564 21184 65570 21248
rect 65254 21183 65570 21184
rect 64334 20704 64650 20705
rect 64334 20640 64340 20704
rect 64404 20640 64420 20704
rect 64484 20640 64500 20704
rect 64564 20640 64580 20704
rect 64644 20640 64650 20704
rect 64334 20639 64650 20640
rect 65254 20160 65570 20161
rect 65254 20096 65260 20160
rect 65324 20096 65340 20160
rect 65404 20096 65420 20160
rect 65484 20096 65500 20160
rect 65564 20096 65570 20160
rect 65254 20095 65570 20096
rect 64334 19616 64650 19617
rect 64334 19552 64340 19616
rect 64404 19552 64420 19616
rect 64484 19552 64500 19616
rect 64564 19552 64580 19616
rect 64644 19552 64650 19616
rect 64334 19551 64650 19552
rect 65254 19072 65570 19073
rect 65254 19008 65260 19072
rect 65324 19008 65340 19072
rect 65404 19008 65420 19072
rect 65484 19008 65500 19072
rect 65564 19008 65570 19072
rect 65254 19007 65570 19008
rect 64334 18528 64650 18529
rect 64334 18464 64340 18528
rect 64404 18464 64420 18528
rect 64484 18464 64500 18528
rect 64564 18464 64580 18528
rect 64644 18464 64650 18528
rect 64334 18463 64650 18464
rect 65254 17984 65570 17985
rect 65254 17920 65260 17984
rect 65324 17920 65340 17984
rect 65404 17920 65420 17984
rect 65484 17920 65500 17984
rect 65564 17920 65570 17984
rect 65254 17919 65570 17920
rect 64334 17440 64650 17441
rect 64334 17376 64340 17440
rect 64404 17376 64420 17440
rect 64484 17376 64500 17440
rect 64564 17376 64580 17440
rect 64644 17376 64650 17440
rect 64334 17375 64650 17376
rect 65254 16896 65570 16897
rect 65254 16832 65260 16896
rect 65324 16832 65340 16896
rect 65404 16832 65420 16896
rect 65484 16832 65500 16896
rect 65564 16832 65570 16896
rect 65254 16831 65570 16832
rect 64965 16690 65031 16693
rect 66069 16690 66135 16693
rect 64965 16688 66135 16690
rect 64965 16632 64970 16688
rect 65026 16632 66074 16688
rect 66130 16632 66135 16688
rect 64965 16630 66135 16632
rect 64965 16627 65031 16630
rect 66069 16627 66135 16630
rect 64334 16352 64650 16353
rect 64334 16288 64340 16352
rect 64404 16288 64420 16352
rect 64484 16288 64500 16352
rect 64564 16288 64580 16352
rect 64644 16288 64650 16352
rect 64334 16287 64650 16288
rect 65254 15808 65570 15809
rect 65254 15744 65260 15808
rect 65324 15744 65340 15808
rect 65404 15744 65420 15808
rect 65484 15744 65500 15808
rect 65564 15744 65570 15808
rect 65254 15743 65570 15744
rect 63350 15268 63356 15332
rect 63420 15330 63426 15332
rect 63420 15270 64154 15330
rect 63420 15268 63426 15270
rect 64094 15197 64154 15270
rect 64334 15264 64650 15265
rect 64334 15200 64340 15264
rect 64404 15200 64420 15264
rect 64484 15200 64500 15264
rect 64564 15200 64580 15264
rect 64644 15200 64650 15264
rect 64334 15199 64650 15200
rect 64094 15192 64203 15197
rect 64094 15136 64142 15192
rect 64198 15136 64203 15192
rect 64094 15134 64203 15136
rect 64137 15131 64203 15134
rect 65254 14720 65570 14721
rect 65254 14656 65260 14720
rect 65324 14656 65340 14720
rect 65404 14656 65420 14720
rect 65484 14656 65500 14720
rect 65564 14656 65570 14720
rect 65254 14655 65570 14656
rect 64334 14176 64650 14177
rect 64334 14112 64340 14176
rect 64404 14112 64420 14176
rect 64484 14112 64500 14176
rect 64564 14112 64580 14176
rect 64644 14112 64650 14176
rect 64334 14111 64650 14112
rect 65254 13632 65570 13633
rect 65254 13568 65260 13632
rect 65324 13568 65340 13632
rect 65404 13568 65420 13632
rect 65484 13568 65500 13632
rect 65564 13568 65570 13632
rect 65254 13567 65570 13568
rect 64334 13088 64650 13089
rect 64334 13024 64340 13088
rect 64404 13024 64420 13088
rect 64484 13024 64500 13088
rect 64564 13024 64580 13088
rect 64644 13024 64650 13088
rect 64334 13023 64650 13024
rect 65254 12544 65570 12545
rect 65254 12480 65260 12544
rect 65324 12480 65340 12544
rect 65404 12480 65420 12544
rect 65484 12480 65500 12544
rect 65564 12480 65570 12544
rect 65254 12479 65570 12480
rect 64334 12000 64650 12001
rect 64334 11936 64340 12000
rect 64404 11936 64420 12000
rect 64484 11936 64500 12000
rect 64564 11936 64580 12000
rect 64644 11936 64650 12000
rect 64334 11935 64650 11936
rect 65254 11456 65570 11457
rect 65254 11392 65260 11456
rect 65324 11392 65340 11456
rect 65404 11392 65420 11456
rect 65484 11392 65500 11456
rect 65564 11392 65570 11456
rect 65254 11391 65570 11392
rect 64334 10912 64650 10913
rect 64334 10848 64340 10912
rect 64404 10848 64420 10912
rect 64484 10848 64500 10912
rect 64564 10848 64580 10912
rect 64644 10848 64650 10912
rect 64334 10847 64650 10848
rect 65254 10368 65570 10369
rect 65254 10304 65260 10368
rect 65324 10304 65340 10368
rect 65404 10304 65420 10368
rect 65484 10304 65500 10368
rect 65564 10304 65570 10368
rect 65254 10303 65570 10304
rect 64334 9824 64650 9825
rect 64334 9760 64340 9824
rect 64404 9760 64420 9824
rect 64484 9760 64500 9824
rect 64564 9760 64580 9824
rect 64644 9760 64650 9824
rect 64334 9759 64650 9760
rect 65254 9280 65570 9281
rect 65254 9216 65260 9280
rect 65324 9216 65340 9280
rect 65404 9216 65420 9280
rect 65484 9216 65500 9280
rect 65564 9216 65570 9280
rect 65254 9215 65570 9216
rect 64334 8736 64650 8737
rect 64334 8672 64340 8736
rect 64404 8672 64420 8736
rect 64484 8672 64500 8736
rect 64564 8672 64580 8736
rect 64644 8672 64650 8736
rect 64334 8671 64650 8672
rect 65254 8192 65570 8193
rect 65254 8128 65260 8192
rect 65324 8128 65340 8192
rect 65404 8128 65420 8192
rect 65484 8128 65500 8192
rect 65564 8128 65570 8192
rect 65254 8127 65570 8128
rect 64334 7648 64650 7649
rect 64334 7584 64340 7648
rect 64404 7584 64420 7648
rect 64484 7584 64500 7648
rect 64564 7584 64580 7648
rect 64644 7584 64650 7648
rect 64334 7583 64650 7584
rect 65254 7104 65570 7105
rect 65254 7040 65260 7104
rect 65324 7040 65340 7104
rect 65404 7040 65420 7104
rect 65484 7040 65500 7104
rect 65564 7040 65570 7104
rect 65254 7039 65570 7040
rect 64334 6560 64650 6561
rect 64334 6496 64340 6560
rect 64404 6496 64420 6560
rect 64484 6496 64500 6560
rect 64564 6496 64580 6560
rect 64644 6496 64650 6560
rect 64334 6495 64650 6496
rect 63902 6020 63908 6084
rect 63972 6082 63978 6084
rect 64689 6082 64755 6085
rect 63972 6080 64755 6082
rect 63972 6024 64694 6080
rect 64750 6024 64755 6080
rect 63972 6022 64755 6024
rect 63972 6020 63978 6022
rect 64689 6019 64755 6022
rect 65254 6016 65570 6017
rect 65254 5952 65260 6016
rect 65324 5952 65340 6016
rect 65404 5952 65420 6016
rect 65484 5952 65500 6016
rect 65564 5952 65570 6016
rect 65254 5951 65570 5952
rect 64137 5948 64203 5949
rect 64086 5884 64092 5948
rect 64156 5946 64203 5948
rect 64156 5944 64248 5946
rect 64198 5888 64248 5944
rect 64156 5886 64248 5888
rect 64156 5884 64203 5886
rect 64137 5883 64203 5884
rect 64334 5472 64650 5473
rect 64334 5408 64340 5472
rect 64404 5408 64420 5472
rect 64484 5408 64500 5472
rect 64564 5408 64580 5472
rect 64644 5408 64650 5472
rect 64334 5407 64650 5408
rect 65254 4928 65570 4929
rect 65254 4864 65260 4928
rect 65324 4864 65340 4928
rect 65404 4864 65420 4928
rect 65484 4864 65500 4928
rect 65564 4864 65570 4928
rect 65254 4863 65570 4864
rect 64334 4384 64650 4385
rect 64334 4320 64340 4384
rect 64404 4320 64420 4384
rect 64484 4320 64500 4384
rect 64564 4320 64580 4384
rect 64644 4320 64650 4384
rect 64334 4319 64650 4320
rect 65254 3840 65570 3841
rect 65254 3776 65260 3840
rect 65324 3776 65340 3840
rect 65404 3776 65420 3840
rect 65484 3776 65500 3840
rect 65564 3776 65570 3840
rect 65254 3775 65570 3776
rect 64334 3296 64650 3297
rect 64334 3232 64340 3296
rect 64404 3232 64420 3296
rect 64484 3232 64500 3296
rect 64564 3232 64580 3296
rect 64644 3232 64650 3296
rect 64334 3231 64650 3232
rect 65254 2752 65570 2753
rect 65254 2688 65260 2752
rect 65324 2688 65340 2752
rect 65404 2688 65420 2752
rect 65484 2688 65500 2752
rect 65564 2688 65570 2752
rect 65254 2687 65570 2688
rect 64334 2208 64650 2209
rect 64334 2144 64340 2208
rect 64404 2144 64420 2208
rect 64484 2144 64500 2208
rect 64564 2144 64580 2208
rect 64644 2144 64650 2208
rect 64334 2143 64650 2144
rect 63718 1940 63724 2004
rect 63788 2002 63794 2004
rect 64689 2002 64755 2005
rect 63788 2000 64755 2002
rect 63788 1944 64694 2000
rect 64750 1944 64755 2000
rect 63788 1942 64755 1944
rect 63788 1940 63794 1942
rect 64689 1939 64755 1942
rect 48957 1868 49023 1869
rect 49233 1868 49299 1869
rect 49693 1868 49759 1869
rect 48935 1866 48941 1868
rect 48866 1806 48941 1866
rect 49005 1864 49023 1868
rect 49211 1866 49217 1868
rect 49018 1808 49023 1864
rect 48935 1804 48941 1806
rect 49005 1804 49023 1808
rect 49142 1806 49217 1866
rect 49281 1864 49299 1868
rect 49668 1866 49674 1868
rect 49294 1808 49299 1864
rect 49211 1804 49217 1806
rect 49281 1804 49299 1808
rect 49602 1806 49674 1866
rect 49738 1864 49759 1868
rect 63493 1866 63559 1869
rect 49754 1808 49759 1864
rect 49668 1804 49674 1806
rect 49738 1804 49759 1808
rect 48957 1803 49023 1804
rect 49233 1803 49299 1804
rect 49693 1803 49759 1804
rect 55170 1864 63559 1866
rect 55170 1808 63498 1864
rect 63554 1808 63559 1864
rect 55170 1806 63559 1808
rect 49366 1668 49372 1732
rect 49436 1730 49442 1732
rect 55170 1730 55230 1806
rect 63493 1803 63559 1806
rect 49436 1670 55230 1730
rect 49436 1668 49442 1670
rect 65254 1664 65570 1665
rect 65254 1600 65260 1664
rect 65324 1600 65340 1664
rect 65404 1600 65420 1664
rect 65484 1600 65500 1664
rect 65564 1600 65570 1664
rect 65254 1599 65570 1600
rect 49073 1532 49079 1596
rect 49143 1594 49149 1596
rect 62849 1594 62915 1597
rect 49143 1592 62915 1594
rect 49143 1536 62854 1592
rect 62910 1536 62915 1592
rect 49143 1534 62915 1536
rect 49143 1532 49149 1534
rect 62849 1531 62915 1534
rect 49918 1260 49924 1324
rect 49988 1322 49994 1324
rect 62573 1322 62639 1325
rect 49988 1320 62639 1322
rect 49988 1264 62578 1320
rect 62634 1264 62639 1320
rect 49988 1262 62639 1264
rect 49988 1260 49994 1262
rect 62573 1259 62639 1262
rect 64334 1120 64650 1121
rect 64334 1056 64340 1120
rect 64404 1056 64420 1120
rect 64484 1056 64500 1120
rect 64564 1056 64580 1120
rect 64644 1056 64650 1120
rect 64334 1055 64650 1056
rect 65254 576 65570 577
rect 65254 512 65260 576
rect 65324 512 65340 576
rect 65404 512 65420 576
rect 65484 512 65500 576
rect 65564 512 65570 576
rect 65254 511 65570 512
<< via3 >>
rect 24348 44916 24412 44980
rect 26004 44916 26068 44980
rect 25452 44780 25516 44844
rect 11652 44644 11716 44708
rect 14964 44644 15028 44708
rect 17724 44644 17788 44708
rect 27660 44644 27724 44708
rect 2000 44636 2064 44640
rect 2000 44580 2004 44636
rect 2004 44580 2060 44636
rect 2060 44580 2064 44636
rect 2000 44576 2064 44580
rect 2080 44636 2144 44640
rect 2080 44580 2084 44636
rect 2084 44580 2140 44636
rect 2140 44580 2144 44636
rect 2080 44576 2144 44580
rect 2160 44636 2224 44640
rect 2160 44580 2164 44636
rect 2164 44580 2220 44636
rect 2220 44580 2224 44636
rect 2160 44576 2224 44580
rect 2240 44636 2304 44640
rect 2240 44580 2244 44636
rect 2244 44580 2300 44636
rect 2300 44580 2304 44636
rect 2240 44576 2304 44580
rect 51000 44636 51064 44640
rect 51000 44580 51004 44636
rect 51004 44580 51060 44636
rect 51060 44580 51064 44636
rect 51000 44576 51064 44580
rect 51080 44636 51144 44640
rect 51080 44580 51084 44636
rect 51084 44580 51140 44636
rect 51140 44580 51144 44636
rect 51080 44576 51144 44580
rect 51160 44636 51224 44640
rect 51160 44580 51164 44636
rect 51164 44580 51220 44636
rect 51220 44580 51224 44636
rect 51160 44576 51224 44580
rect 51240 44636 51304 44640
rect 51240 44580 51244 44636
rect 51244 44580 51300 44636
rect 51300 44580 51304 44636
rect 51240 44576 51304 44580
rect 6132 44568 6196 44572
rect 6132 44512 6182 44568
rect 6182 44512 6196 44568
rect 6132 44508 6196 44512
rect 6684 44568 6748 44572
rect 6684 44512 6734 44568
rect 6734 44512 6748 44568
rect 6684 44508 6748 44512
rect 7236 44568 7300 44572
rect 7236 44512 7286 44568
rect 7286 44512 7300 44568
rect 7236 44508 7300 44512
rect 7788 44568 7852 44572
rect 7788 44512 7838 44568
rect 7838 44512 7852 44568
rect 7788 44508 7852 44512
rect 8340 44568 8404 44572
rect 8340 44512 8390 44568
rect 8390 44512 8404 44568
rect 8340 44508 8404 44512
rect 8892 44568 8956 44572
rect 8892 44512 8942 44568
rect 8942 44512 8956 44568
rect 8892 44508 8956 44512
rect 9444 44568 9508 44572
rect 9444 44512 9494 44568
rect 9494 44512 9508 44568
rect 9444 44508 9508 44512
rect 9996 44568 10060 44572
rect 9996 44512 10046 44568
rect 10046 44512 10060 44568
rect 9996 44508 10060 44512
rect 10548 44568 10612 44572
rect 10548 44512 10598 44568
rect 10598 44512 10612 44568
rect 10548 44508 10612 44512
rect 12204 44568 12268 44572
rect 12204 44512 12254 44568
rect 12254 44512 12268 44568
rect 12204 44508 12268 44512
rect 12756 44568 12820 44572
rect 12756 44512 12806 44568
rect 12806 44512 12820 44568
rect 12756 44508 12820 44512
rect 13308 44508 13372 44572
rect 13860 44568 13924 44572
rect 13860 44512 13874 44568
rect 13874 44512 13924 44568
rect 13860 44508 13924 44512
rect 15516 44568 15580 44572
rect 15516 44512 15530 44568
rect 15530 44512 15580 44568
rect 15516 44508 15580 44512
rect 16068 44508 16132 44572
rect 16620 44568 16684 44572
rect 16620 44512 16670 44568
rect 16670 44512 16684 44568
rect 16620 44508 16684 44512
rect 17172 44508 17236 44572
rect 26556 44372 26620 44436
rect 27108 44372 27172 44436
rect 28212 44372 28276 44436
rect 2920 44092 2984 44096
rect 2920 44036 2924 44092
rect 2924 44036 2980 44092
rect 2980 44036 2984 44092
rect 2920 44032 2984 44036
rect 3000 44092 3064 44096
rect 3000 44036 3004 44092
rect 3004 44036 3060 44092
rect 3060 44036 3064 44092
rect 3000 44032 3064 44036
rect 3080 44092 3144 44096
rect 3080 44036 3084 44092
rect 3084 44036 3140 44092
rect 3140 44036 3144 44092
rect 3080 44032 3144 44036
rect 3160 44092 3224 44096
rect 3160 44036 3164 44092
rect 3164 44036 3220 44092
rect 3220 44036 3224 44092
rect 3160 44032 3224 44036
rect 51920 44092 51984 44096
rect 51920 44036 51924 44092
rect 51924 44036 51980 44092
rect 51980 44036 51984 44092
rect 51920 44032 51984 44036
rect 52000 44092 52064 44096
rect 52000 44036 52004 44092
rect 52004 44036 52060 44092
rect 52060 44036 52064 44092
rect 52000 44032 52064 44036
rect 52080 44092 52144 44096
rect 52080 44036 52084 44092
rect 52084 44036 52140 44092
rect 52140 44036 52144 44092
rect 52080 44032 52144 44036
rect 52160 44092 52224 44096
rect 52160 44036 52164 44092
rect 52164 44036 52220 44092
rect 52220 44036 52224 44092
rect 52160 44032 52224 44036
rect 11100 43888 11164 43892
rect 11100 43832 11150 43888
rect 11150 43832 11164 43888
rect 11100 43828 11164 43832
rect 14412 43828 14476 43892
rect 18828 43692 18892 43756
rect 31892 43692 31956 43756
rect 2000 43548 2064 43552
rect 2000 43492 2004 43548
rect 2004 43492 2060 43548
rect 2060 43492 2064 43548
rect 2000 43488 2064 43492
rect 2080 43548 2144 43552
rect 2080 43492 2084 43548
rect 2084 43492 2140 43548
rect 2140 43492 2144 43548
rect 2080 43488 2144 43492
rect 2160 43548 2224 43552
rect 2160 43492 2164 43548
rect 2164 43492 2220 43548
rect 2220 43492 2224 43548
rect 2160 43488 2224 43492
rect 2240 43548 2304 43552
rect 2240 43492 2244 43548
rect 2244 43492 2300 43548
rect 2300 43492 2304 43548
rect 2240 43488 2304 43492
rect 51000 43548 51064 43552
rect 51000 43492 51004 43548
rect 51004 43492 51060 43548
rect 51060 43492 51064 43548
rect 51000 43488 51064 43492
rect 51080 43548 51144 43552
rect 51080 43492 51084 43548
rect 51084 43492 51140 43548
rect 51140 43492 51144 43548
rect 51080 43488 51144 43492
rect 51160 43548 51224 43552
rect 51160 43492 51164 43548
rect 51164 43492 51220 43548
rect 51220 43492 51224 43548
rect 51160 43488 51224 43492
rect 51240 43548 51304 43552
rect 51240 43492 51244 43548
rect 51244 43492 51300 43548
rect 51300 43492 51304 43548
rect 51240 43488 51304 43492
rect 18276 43420 18340 43484
rect 22692 43148 22756 43212
rect 24532 43148 24596 43212
rect 27108 43012 27172 43076
rect 2920 43004 2984 43008
rect 2920 42948 2924 43004
rect 2924 42948 2980 43004
rect 2980 42948 2984 43004
rect 2920 42944 2984 42948
rect 3000 43004 3064 43008
rect 3000 42948 3004 43004
rect 3004 42948 3060 43004
rect 3060 42948 3064 43004
rect 3000 42944 3064 42948
rect 3080 43004 3144 43008
rect 3080 42948 3084 43004
rect 3084 42948 3140 43004
rect 3140 42948 3144 43004
rect 3080 42944 3144 42948
rect 3160 43004 3224 43008
rect 3160 42948 3164 43004
rect 3164 42948 3220 43004
rect 3220 42948 3224 43004
rect 3160 42944 3224 42948
rect 51920 43004 51984 43008
rect 51920 42948 51924 43004
rect 51924 42948 51980 43004
rect 51980 42948 51984 43004
rect 51920 42944 51984 42948
rect 52000 43004 52064 43008
rect 52000 42948 52004 43004
rect 52004 42948 52060 43004
rect 52060 42948 52064 43004
rect 52000 42944 52064 42948
rect 52080 43004 52144 43008
rect 52080 42948 52084 43004
rect 52084 42948 52140 43004
rect 52140 42948 52144 43004
rect 52080 42944 52144 42948
rect 52160 43004 52224 43008
rect 52160 42948 52164 43004
rect 52164 42948 52220 43004
rect 52220 42948 52224 43004
rect 52160 42944 52224 42948
rect 23244 42740 23308 42804
rect 28948 42740 29012 42804
rect 2000 42460 2064 42464
rect 2000 42404 2004 42460
rect 2004 42404 2060 42460
rect 2060 42404 2064 42460
rect 2000 42400 2064 42404
rect 2080 42460 2144 42464
rect 2080 42404 2084 42460
rect 2084 42404 2140 42460
rect 2140 42404 2144 42460
rect 2080 42400 2144 42404
rect 2160 42460 2224 42464
rect 2160 42404 2164 42460
rect 2164 42404 2220 42460
rect 2220 42404 2224 42460
rect 2160 42400 2224 42404
rect 2240 42460 2304 42464
rect 2240 42404 2244 42460
rect 2244 42404 2300 42460
rect 2300 42404 2304 42460
rect 2240 42400 2304 42404
rect 51000 42460 51064 42464
rect 51000 42404 51004 42460
rect 51004 42404 51060 42460
rect 51060 42404 51064 42460
rect 51000 42400 51064 42404
rect 51080 42460 51144 42464
rect 51080 42404 51084 42460
rect 51084 42404 51140 42460
rect 51140 42404 51144 42460
rect 51080 42400 51144 42404
rect 51160 42460 51224 42464
rect 51160 42404 51164 42460
rect 51164 42404 51220 42460
rect 51220 42404 51224 42460
rect 51160 42400 51224 42404
rect 51240 42460 51304 42464
rect 51240 42404 51244 42460
rect 51244 42404 51300 42460
rect 51300 42404 51304 42460
rect 51240 42400 51304 42404
rect 27844 42332 27908 42396
rect 28212 42196 28276 42260
rect 62620 42196 62684 42260
rect 17908 42060 17972 42124
rect 30972 41924 31036 41988
rect 2920 41916 2984 41920
rect 2920 41860 2924 41916
rect 2924 41860 2980 41916
rect 2980 41860 2984 41916
rect 2920 41856 2984 41860
rect 3000 41916 3064 41920
rect 3000 41860 3004 41916
rect 3004 41860 3060 41916
rect 3060 41860 3064 41916
rect 3000 41856 3064 41860
rect 3080 41916 3144 41920
rect 3080 41860 3084 41916
rect 3084 41860 3140 41916
rect 3140 41860 3144 41916
rect 3080 41856 3144 41860
rect 3160 41916 3224 41920
rect 3160 41860 3164 41916
rect 3164 41860 3220 41916
rect 3220 41860 3224 41916
rect 3160 41856 3224 41860
rect 51920 41916 51984 41920
rect 51920 41860 51924 41916
rect 51924 41860 51980 41916
rect 51980 41860 51984 41916
rect 51920 41856 51984 41860
rect 52000 41916 52064 41920
rect 52000 41860 52004 41916
rect 52004 41860 52060 41916
rect 52060 41860 52064 41916
rect 52000 41856 52064 41860
rect 52080 41916 52144 41920
rect 52080 41860 52084 41916
rect 52084 41860 52140 41916
rect 52140 41860 52144 41916
rect 52080 41856 52144 41860
rect 52160 41916 52224 41920
rect 52160 41860 52164 41916
rect 52164 41860 52220 41916
rect 52220 41860 52224 41916
rect 52160 41856 52224 41860
rect 36124 41652 36188 41716
rect 35020 41380 35084 41444
rect 2000 41372 2064 41376
rect 2000 41316 2004 41372
rect 2004 41316 2060 41372
rect 2060 41316 2064 41372
rect 2000 41312 2064 41316
rect 2080 41372 2144 41376
rect 2080 41316 2084 41372
rect 2084 41316 2140 41372
rect 2140 41316 2144 41372
rect 2080 41312 2144 41316
rect 2160 41372 2224 41376
rect 2160 41316 2164 41372
rect 2164 41316 2220 41372
rect 2220 41316 2224 41372
rect 2160 41312 2224 41316
rect 2240 41372 2304 41376
rect 2240 41316 2244 41372
rect 2244 41316 2300 41372
rect 2300 41316 2304 41372
rect 2240 41312 2304 41316
rect 51000 41372 51064 41376
rect 51000 41316 51004 41372
rect 51004 41316 51060 41372
rect 51060 41316 51064 41372
rect 51000 41312 51064 41316
rect 51080 41372 51144 41376
rect 51080 41316 51084 41372
rect 51084 41316 51140 41372
rect 51140 41316 51144 41372
rect 51080 41312 51144 41316
rect 51160 41372 51224 41376
rect 51160 41316 51164 41372
rect 51164 41316 51220 41372
rect 51220 41316 51224 41372
rect 51160 41312 51224 41316
rect 51240 41372 51304 41376
rect 51240 41316 51244 41372
rect 51244 41316 51300 41372
rect 51300 41316 51304 41372
rect 51240 41312 51304 41316
rect 26740 41244 26804 41308
rect 22140 41108 22204 41172
rect 28948 40972 29012 41036
rect 32996 40836 33060 40900
rect 2920 40828 2984 40832
rect 2920 40772 2924 40828
rect 2924 40772 2980 40828
rect 2980 40772 2984 40828
rect 2920 40768 2984 40772
rect 3000 40828 3064 40832
rect 3000 40772 3004 40828
rect 3004 40772 3060 40828
rect 3060 40772 3064 40828
rect 3000 40768 3064 40772
rect 3080 40828 3144 40832
rect 3080 40772 3084 40828
rect 3084 40772 3140 40828
rect 3140 40772 3144 40828
rect 3080 40768 3144 40772
rect 3160 40828 3224 40832
rect 3160 40772 3164 40828
rect 3164 40772 3220 40828
rect 3220 40772 3224 40828
rect 3160 40768 3224 40772
rect 51920 40828 51984 40832
rect 51920 40772 51924 40828
rect 51924 40772 51980 40828
rect 51980 40772 51984 40828
rect 51920 40768 51984 40772
rect 52000 40828 52064 40832
rect 52000 40772 52004 40828
rect 52004 40772 52060 40828
rect 52060 40772 52064 40828
rect 52000 40768 52064 40772
rect 52080 40828 52144 40832
rect 52080 40772 52084 40828
rect 52084 40772 52140 40828
rect 52140 40772 52144 40828
rect 52080 40768 52144 40772
rect 52160 40828 52224 40832
rect 52160 40772 52164 40828
rect 52164 40772 52220 40828
rect 52220 40772 52224 40828
rect 52160 40768 52224 40772
rect 2000 40284 2064 40288
rect 2000 40228 2004 40284
rect 2004 40228 2060 40284
rect 2060 40228 2064 40284
rect 2000 40224 2064 40228
rect 2080 40284 2144 40288
rect 2080 40228 2084 40284
rect 2084 40228 2140 40284
rect 2140 40228 2144 40284
rect 2080 40224 2144 40228
rect 2160 40284 2224 40288
rect 2160 40228 2164 40284
rect 2164 40228 2220 40284
rect 2220 40228 2224 40284
rect 2160 40224 2224 40228
rect 2240 40284 2304 40288
rect 2240 40228 2244 40284
rect 2244 40228 2300 40284
rect 2300 40228 2304 40284
rect 2240 40224 2304 40228
rect 51000 40284 51064 40288
rect 51000 40228 51004 40284
rect 51004 40228 51060 40284
rect 51060 40228 51064 40284
rect 51000 40224 51064 40228
rect 51080 40284 51144 40288
rect 51080 40228 51084 40284
rect 51084 40228 51140 40284
rect 51140 40228 51144 40284
rect 51080 40224 51144 40228
rect 51160 40284 51224 40288
rect 51160 40228 51164 40284
rect 51164 40228 51220 40284
rect 51220 40228 51224 40284
rect 51160 40224 51224 40228
rect 51240 40284 51304 40288
rect 51240 40228 51244 40284
rect 51244 40228 51300 40284
rect 51300 40228 51304 40284
rect 51240 40224 51304 40228
rect 32076 40080 32140 40084
rect 44588 40156 44652 40220
rect 63540 40156 63604 40220
rect 32076 40024 32090 40080
rect 32090 40024 32140 40080
rect 32076 40020 32140 40024
rect 19012 39748 19076 39812
rect 2920 39740 2984 39744
rect 2920 39684 2924 39740
rect 2924 39684 2980 39740
rect 2980 39684 2984 39740
rect 2920 39680 2984 39684
rect 3000 39740 3064 39744
rect 3000 39684 3004 39740
rect 3004 39684 3060 39740
rect 3060 39684 3064 39740
rect 3000 39680 3064 39684
rect 3080 39740 3144 39744
rect 3080 39684 3084 39740
rect 3084 39684 3140 39740
rect 3140 39684 3144 39740
rect 3080 39680 3144 39684
rect 3160 39740 3224 39744
rect 3160 39684 3164 39740
rect 3164 39684 3220 39740
rect 3220 39684 3224 39740
rect 3160 39680 3224 39684
rect 31892 39748 31956 39812
rect 46980 39748 47044 39812
rect 51920 39740 51984 39744
rect 51920 39684 51924 39740
rect 51924 39684 51980 39740
rect 51980 39684 51984 39740
rect 51920 39680 51984 39684
rect 52000 39740 52064 39744
rect 52000 39684 52004 39740
rect 52004 39684 52060 39740
rect 52060 39684 52064 39740
rect 52000 39680 52064 39684
rect 52080 39740 52144 39744
rect 52080 39684 52084 39740
rect 52084 39684 52140 39740
rect 52140 39684 52144 39740
rect 52080 39680 52144 39684
rect 52160 39740 52224 39744
rect 52160 39684 52164 39740
rect 52164 39684 52220 39740
rect 52220 39684 52224 39740
rect 52160 39680 52224 39684
rect 26004 39476 26068 39540
rect 31340 39476 31404 39540
rect 15516 39340 15580 39404
rect 28948 39340 29012 39404
rect 22508 39204 22572 39268
rect 2000 39196 2064 39200
rect 2000 39140 2004 39196
rect 2004 39140 2060 39196
rect 2060 39140 2064 39196
rect 2000 39136 2064 39140
rect 2080 39196 2144 39200
rect 2080 39140 2084 39196
rect 2084 39140 2140 39196
rect 2140 39140 2144 39196
rect 2080 39136 2144 39140
rect 2160 39196 2224 39200
rect 2160 39140 2164 39196
rect 2164 39140 2220 39196
rect 2220 39140 2224 39196
rect 2160 39136 2224 39140
rect 2240 39196 2304 39200
rect 2240 39140 2244 39196
rect 2244 39140 2300 39196
rect 2300 39140 2304 39196
rect 2240 39136 2304 39140
rect 51000 39196 51064 39200
rect 51000 39140 51004 39196
rect 51004 39140 51060 39196
rect 51060 39140 51064 39196
rect 51000 39136 51064 39140
rect 51080 39196 51144 39200
rect 51080 39140 51084 39196
rect 51084 39140 51140 39196
rect 51140 39140 51144 39196
rect 51080 39136 51144 39140
rect 51160 39196 51224 39200
rect 51160 39140 51164 39196
rect 51164 39140 51220 39196
rect 51220 39140 51224 39196
rect 51160 39136 51224 39140
rect 51240 39196 51304 39200
rect 51240 39140 51244 39196
rect 51244 39140 51300 39196
rect 51300 39140 51304 39196
rect 51240 39136 51304 39140
rect 27292 39068 27356 39132
rect 24532 38796 24596 38860
rect 27476 38796 27540 38860
rect 28396 38660 28460 38724
rect 2920 38652 2984 38656
rect 2920 38596 2924 38652
rect 2924 38596 2980 38652
rect 2980 38596 2984 38652
rect 2920 38592 2984 38596
rect 3000 38652 3064 38656
rect 3000 38596 3004 38652
rect 3004 38596 3060 38652
rect 3060 38596 3064 38652
rect 3000 38592 3064 38596
rect 3080 38652 3144 38656
rect 3080 38596 3084 38652
rect 3084 38596 3140 38652
rect 3140 38596 3144 38652
rect 3080 38592 3144 38596
rect 3160 38652 3224 38656
rect 3160 38596 3164 38652
rect 3164 38596 3220 38652
rect 3220 38596 3224 38652
rect 3160 38592 3224 38596
rect 51920 38652 51984 38656
rect 51920 38596 51924 38652
rect 51924 38596 51980 38652
rect 51980 38596 51984 38652
rect 51920 38592 51984 38596
rect 52000 38652 52064 38656
rect 52000 38596 52004 38652
rect 52004 38596 52060 38652
rect 52060 38596 52064 38652
rect 52000 38592 52064 38596
rect 52080 38652 52144 38656
rect 52080 38596 52084 38652
rect 52084 38596 52140 38652
rect 52140 38596 52144 38652
rect 52080 38592 52144 38596
rect 52160 38652 52224 38656
rect 52160 38596 52164 38652
rect 52164 38596 52220 38652
rect 52220 38596 52224 38652
rect 52160 38592 52224 38596
rect 35388 38524 35452 38588
rect 21404 38252 21468 38316
rect 32996 38252 33060 38316
rect 2000 38108 2064 38112
rect 2000 38052 2004 38108
rect 2004 38052 2060 38108
rect 2060 38052 2064 38108
rect 2000 38048 2064 38052
rect 2080 38108 2144 38112
rect 2080 38052 2084 38108
rect 2084 38052 2140 38108
rect 2140 38052 2144 38108
rect 2080 38048 2144 38052
rect 2160 38108 2224 38112
rect 2160 38052 2164 38108
rect 2164 38052 2220 38108
rect 2220 38052 2224 38108
rect 2160 38048 2224 38052
rect 2240 38108 2304 38112
rect 2240 38052 2244 38108
rect 2244 38052 2300 38108
rect 2300 38052 2304 38108
rect 2240 38048 2304 38052
rect 14412 37980 14476 38044
rect 51000 38108 51064 38112
rect 51000 38052 51004 38108
rect 51004 38052 51060 38108
rect 51060 38052 51064 38108
rect 51000 38048 51064 38052
rect 51080 38108 51144 38112
rect 51080 38052 51084 38108
rect 51084 38052 51140 38108
rect 51140 38052 51144 38108
rect 51080 38048 51144 38052
rect 51160 38108 51224 38112
rect 51160 38052 51164 38108
rect 51164 38052 51220 38108
rect 51220 38052 51224 38108
rect 51160 38048 51224 38052
rect 51240 38108 51304 38112
rect 51240 38052 51244 38108
rect 51244 38052 51300 38108
rect 51300 38052 51304 38108
rect 51240 38048 51304 38052
rect 24900 37980 24964 38044
rect 27476 37844 27540 37908
rect 30236 37844 30300 37908
rect 32076 37844 32140 37908
rect 32996 37844 33060 37908
rect 20116 37572 20180 37636
rect 2920 37564 2984 37568
rect 2920 37508 2924 37564
rect 2924 37508 2980 37564
rect 2980 37508 2984 37564
rect 2920 37504 2984 37508
rect 3000 37564 3064 37568
rect 3000 37508 3004 37564
rect 3004 37508 3060 37564
rect 3060 37508 3064 37564
rect 3000 37504 3064 37508
rect 3080 37564 3144 37568
rect 3080 37508 3084 37564
rect 3084 37508 3140 37564
rect 3140 37508 3144 37564
rect 3080 37504 3144 37508
rect 3160 37564 3224 37568
rect 3160 37508 3164 37564
rect 3164 37508 3220 37564
rect 3220 37508 3224 37564
rect 3160 37504 3224 37508
rect 51920 37564 51984 37568
rect 51920 37508 51924 37564
rect 51924 37508 51980 37564
rect 51980 37508 51984 37564
rect 51920 37504 51984 37508
rect 52000 37564 52064 37568
rect 52000 37508 52004 37564
rect 52004 37508 52060 37564
rect 52060 37508 52064 37564
rect 52000 37504 52064 37508
rect 52080 37564 52144 37568
rect 52080 37508 52084 37564
rect 52084 37508 52140 37564
rect 52140 37508 52144 37564
rect 52080 37504 52144 37508
rect 52160 37564 52224 37568
rect 52160 37508 52164 37564
rect 52164 37508 52220 37564
rect 52220 37508 52224 37564
rect 52160 37504 52224 37508
rect 65260 37564 65324 37568
rect 65260 37508 65264 37564
rect 65264 37508 65320 37564
rect 65320 37508 65324 37564
rect 65260 37504 65324 37508
rect 65340 37564 65404 37568
rect 65340 37508 65344 37564
rect 65344 37508 65400 37564
rect 65400 37508 65404 37564
rect 65340 37504 65404 37508
rect 65420 37564 65484 37568
rect 65420 37508 65424 37564
rect 65424 37508 65480 37564
rect 65480 37508 65484 37564
rect 65420 37504 65484 37508
rect 65500 37564 65564 37568
rect 65500 37508 65504 37564
rect 65504 37508 65560 37564
rect 65560 37508 65564 37564
rect 65500 37504 65564 37508
rect 29316 37436 29380 37500
rect 32076 37300 32140 37364
rect 32444 37224 32508 37228
rect 33732 37360 33796 37364
rect 33732 37304 33746 37360
rect 33746 37304 33796 37360
rect 33732 37300 33796 37304
rect 32444 37168 32458 37224
rect 32458 37168 32508 37224
rect 32444 37164 32508 37168
rect 33364 37164 33428 37228
rect 42380 37164 42444 37228
rect 10916 37028 10980 37092
rect 21036 37028 21100 37092
rect 32812 37028 32876 37092
rect 2000 37020 2064 37024
rect 2000 36964 2004 37020
rect 2004 36964 2060 37020
rect 2060 36964 2064 37020
rect 2000 36960 2064 36964
rect 2080 37020 2144 37024
rect 2080 36964 2084 37020
rect 2084 36964 2140 37020
rect 2140 36964 2144 37020
rect 2080 36960 2144 36964
rect 2160 37020 2224 37024
rect 2160 36964 2164 37020
rect 2164 36964 2220 37020
rect 2220 36964 2224 37020
rect 2160 36960 2224 36964
rect 2240 37020 2304 37024
rect 2240 36964 2244 37020
rect 2244 36964 2300 37020
rect 2300 36964 2304 37020
rect 2240 36960 2304 36964
rect 51000 37020 51064 37024
rect 51000 36964 51004 37020
rect 51004 36964 51060 37020
rect 51060 36964 51064 37020
rect 51000 36960 51064 36964
rect 51080 37020 51144 37024
rect 51080 36964 51084 37020
rect 51084 36964 51140 37020
rect 51140 36964 51144 37020
rect 51080 36960 51144 36964
rect 51160 37020 51224 37024
rect 51160 36964 51164 37020
rect 51164 36964 51220 37020
rect 51220 36964 51224 37020
rect 51160 36960 51224 36964
rect 51240 37020 51304 37024
rect 51240 36964 51244 37020
rect 51244 36964 51300 37020
rect 51300 36964 51304 37020
rect 51240 36960 51304 36964
rect 64340 37020 64404 37024
rect 64340 36964 64344 37020
rect 64344 36964 64400 37020
rect 64400 36964 64404 37020
rect 64340 36960 64404 36964
rect 64420 37020 64484 37024
rect 64420 36964 64424 37020
rect 64424 36964 64480 37020
rect 64480 36964 64484 37020
rect 64420 36960 64484 36964
rect 64500 37020 64564 37024
rect 64500 36964 64504 37020
rect 64504 36964 64560 37020
rect 64560 36964 64564 37020
rect 64500 36960 64564 36964
rect 64580 37020 64644 37024
rect 64580 36964 64584 37020
rect 64584 36964 64640 37020
rect 64640 36964 64644 37020
rect 64580 36960 64644 36964
rect 9628 36892 9692 36956
rect 21588 36952 21652 36956
rect 21588 36896 21638 36952
rect 21638 36896 21652 36952
rect 21588 36892 21652 36896
rect 23796 36892 23860 36956
rect 12020 36756 12084 36820
rect 30604 36756 30668 36820
rect 45876 36756 45940 36820
rect 6132 36620 6196 36684
rect 39988 36620 40052 36684
rect 3924 36484 3988 36548
rect 23612 36484 23676 36548
rect 65260 36476 65324 36480
rect 65260 36420 65264 36476
rect 65264 36420 65320 36476
rect 65320 36420 65324 36476
rect 65260 36416 65324 36420
rect 65340 36476 65404 36480
rect 65340 36420 65344 36476
rect 65344 36420 65400 36476
rect 65400 36420 65404 36476
rect 65340 36416 65404 36420
rect 65420 36476 65484 36480
rect 65420 36420 65424 36476
rect 65424 36420 65480 36476
rect 65480 36420 65484 36476
rect 65420 36416 65484 36420
rect 65500 36476 65564 36480
rect 65500 36420 65504 36476
rect 65504 36420 65560 36476
rect 65560 36420 65564 36476
rect 65500 36416 65564 36420
rect 25084 36348 25148 36412
rect 64092 36348 64156 36412
rect 19564 36212 19628 36276
rect 16620 36076 16684 36140
rect 4982 35940 5046 36004
rect 13158 35940 13222 36004
rect 26474 35940 26538 36004
rect 34044 35940 34108 36004
rect 63908 36212 63972 36276
rect 37686 35940 37750 36004
rect 63356 35940 63420 36004
rect 64340 35932 64404 35936
rect 64340 35876 64344 35932
rect 64344 35876 64400 35932
rect 64400 35876 64404 35932
rect 64340 35872 64404 35876
rect 64420 35932 64484 35936
rect 64420 35876 64424 35932
rect 64424 35876 64480 35932
rect 64480 35876 64484 35932
rect 64420 35872 64484 35876
rect 64500 35932 64564 35936
rect 64500 35876 64504 35932
rect 64504 35876 64560 35932
rect 64560 35876 64564 35932
rect 64500 35872 64564 35876
rect 64580 35932 64644 35936
rect 64580 35876 64584 35932
rect 64584 35876 64640 35932
rect 64640 35876 64644 35932
rect 64580 35872 64644 35876
rect 21968 35864 22032 35868
rect 21968 35808 22006 35864
rect 22006 35808 22032 35864
rect 21968 35804 22032 35808
rect 23532 35864 23596 35868
rect 23532 35808 23570 35864
rect 23570 35808 23596 35864
rect 23532 35804 23596 35808
rect 24474 35864 24538 35868
rect 24474 35808 24490 35864
rect 24490 35808 24538 35864
rect 24474 35804 24538 35808
rect 24716 35864 24780 35868
rect 24716 35808 24766 35864
rect 24766 35808 24780 35864
rect 24716 35804 24780 35808
rect 25868 35864 25932 35868
rect 25868 35808 25870 35864
rect 25870 35808 25926 35864
rect 25926 35808 25932 35864
rect 25868 35804 25932 35808
rect 29510 35804 29574 35868
rect 30198 35864 30262 35868
rect 30198 35808 30250 35864
rect 30250 35808 30262 35864
rect 30198 35804 30262 35808
rect 30696 35804 30760 35868
rect 7328 35668 7392 35732
rect 8486 35668 8550 35732
rect 20028 35728 20092 35732
rect 20028 35672 20074 35728
rect 20074 35672 20092 35728
rect 20028 35668 20092 35672
rect 21196 35668 21260 35732
rect 22198 35728 22262 35732
rect 22198 35672 22246 35728
rect 22246 35672 22262 35728
rect 22198 35668 22262 35672
rect 22968 35728 23032 35732
rect 22968 35672 23018 35728
rect 23018 35672 23032 35728
rect 22968 35668 23032 35672
rect 23198 35728 23262 35732
rect 23198 35672 23202 35728
rect 23202 35672 23258 35728
rect 23258 35672 23262 35728
rect 23198 35668 23262 35672
rect 25210 35728 25274 35732
rect 25210 35672 25226 35728
rect 25226 35672 25274 35728
rect 25210 35668 25274 35672
rect 29968 35668 30032 35732
rect 31846 35804 31910 35868
rect 34182 35804 34246 35868
rect 35198 35804 35262 35868
rect 38854 35804 38918 35868
rect 43526 35804 43590 35868
rect 36518 35728 36582 35732
rect 36518 35672 36542 35728
rect 36542 35672 36582 35728
rect 36518 35668 36582 35672
rect 41184 35668 41248 35732
rect 56246 35668 56310 35732
rect 2000 35428 2064 35492
rect 2080 35428 2144 35492
rect 2160 35428 2224 35492
rect 2240 35428 2304 35492
rect 2000 35348 2064 35412
rect 2080 35348 2144 35412
rect 2160 35348 2224 35412
rect 2240 35348 2304 35412
rect 2000 35268 2064 35332
rect 2080 35268 2144 35332
rect 2160 35268 2224 35332
rect 2240 35268 2304 35332
rect 2000 35188 2064 35252
rect 2080 35188 2144 35252
rect 2160 35188 2224 35252
rect 2240 35188 2304 35252
rect 51000 35428 51064 35492
rect 51080 35428 51144 35492
rect 51160 35428 51224 35492
rect 51240 35428 51304 35492
rect 51000 35348 51064 35412
rect 51080 35348 51144 35412
rect 51160 35348 51224 35412
rect 51240 35348 51304 35412
rect 51000 35268 51064 35332
rect 51080 35268 51144 35332
rect 51160 35268 51224 35332
rect 51240 35268 51304 35332
rect 65260 35388 65324 35392
rect 65260 35332 65264 35388
rect 65264 35332 65320 35388
rect 65320 35332 65324 35388
rect 65260 35328 65324 35332
rect 65340 35388 65404 35392
rect 65340 35332 65344 35388
rect 65344 35332 65400 35388
rect 65400 35332 65404 35388
rect 65340 35328 65404 35332
rect 65420 35388 65484 35392
rect 65420 35332 65424 35388
rect 65424 35332 65480 35388
rect 65480 35332 65484 35388
rect 65420 35328 65484 35332
rect 65500 35388 65564 35392
rect 65500 35332 65504 35388
rect 65504 35332 65560 35388
rect 65560 35332 65564 35388
rect 65500 35328 65564 35332
rect 51000 35188 51064 35252
rect 51080 35188 51144 35252
rect 51160 35188 51224 35252
rect 51240 35188 51304 35252
rect 2920 34732 2984 34796
rect 3000 34732 3064 34796
rect 3080 34732 3144 34796
rect 3160 34732 3224 34796
rect 2920 34652 2984 34716
rect 3000 34652 3064 34716
rect 3080 34652 3144 34716
rect 3160 34652 3224 34716
rect 2920 34572 2984 34636
rect 3000 34572 3064 34636
rect 3080 34572 3144 34636
rect 3160 34572 3224 34636
rect 2920 34492 2984 34556
rect 3000 34492 3064 34556
rect 3080 34492 3144 34556
rect 3160 34492 3224 34556
rect 51920 34732 51984 34796
rect 52000 34732 52064 34796
rect 52080 34732 52144 34796
rect 52160 34732 52224 34796
rect 64340 34844 64404 34848
rect 64340 34788 64344 34844
rect 64344 34788 64400 34844
rect 64400 34788 64404 34844
rect 64340 34784 64404 34788
rect 64420 34844 64484 34848
rect 64420 34788 64424 34844
rect 64424 34788 64480 34844
rect 64480 34788 64484 34844
rect 64420 34784 64484 34788
rect 64500 34844 64564 34848
rect 64500 34788 64504 34844
rect 64504 34788 64560 34844
rect 64560 34788 64564 34844
rect 64500 34784 64564 34788
rect 64580 34844 64644 34848
rect 64580 34788 64584 34844
rect 64584 34788 64640 34844
rect 64640 34788 64644 34844
rect 64580 34784 64644 34788
rect 51920 34652 51984 34716
rect 52000 34652 52064 34716
rect 52080 34652 52144 34716
rect 52160 34652 52224 34716
rect 63724 34716 63788 34780
rect 51920 34572 51984 34636
rect 52000 34572 52064 34636
rect 52080 34572 52144 34636
rect 52160 34572 52224 34636
rect 63540 34580 63604 34644
rect 51920 34492 51984 34556
rect 52000 34492 52064 34556
rect 52080 34492 52144 34556
rect 52160 34492 52224 34556
rect 65260 34300 65324 34304
rect 65260 34244 65264 34300
rect 65264 34244 65320 34300
rect 65320 34244 65324 34300
rect 65260 34240 65324 34244
rect 65340 34300 65404 34304
rect 65340 34244 65344 34300
rect 65344 34244 65400 34300
rect 65400 34244 65404 34300
rect 65340 34240 65404 34244
rect 65420 34300 65484 34304
rect 65420 34244 65424 34300
rect 65424 34244 65480 34300
rect 65480 34244 65484 34300
rect 65420 34240 65484 34244
rect 65500 34300 65564 34304
rect 65500 34244 65504 34300
rect 65504 34244 65560 34300
rect 65560 34244 65564 34300
rect 65500 34240 65564 34244
rect 64340 33756 64404 33760
rect 64340 33700 64344 33756
rect 64344 33700 64400 33756
rect 64400 33700 64404 33756
rect 64340 33696 64404 33700
rect 64420 33756 64484 33760
rect 64420 33700 64424 33756
rect 64424 33700 64480 33756
rect 64480 33700 64484 33756
rect 64420 33696 64484 33700
rect 64500 33756 64564 33760
rect 64500 33700 64504 33756
rect 64504 33700 64560 33756
rect 64560 33700 64564 33756
rect 64500 33696 64564 33700
rect 64580 33756 64644 33760
rect 64580 33700 64584 33756
rect 64584 33700 64640 33756
rect 64640 33700 64644 33756
rect 64580 33696 64644 33700
rect 65260 33212 65324 33216
rect 65260 33156 65264 33212
rect 65264 33156 65320 33212
rect 65320 33156 65324 33212
rect 65260 33152 65324 33156
rect 65340 33212 65404 33216
rect 65340 33156 65344 33212
rect 65344 33156 65400 33212
rect 65400 33156 65404 33212
rect 65340 33152 65404 33156
rect 65420 33212 65484 33216
rect 65420 33156 65424 33212
rect 65424 33156 65480 33212
rect 65480 33156 65484 33212
rect 65420 33152 65484 33156
rect 65500 33212 65564 33216
rect 65500 33156 65504 33212
rect 65504 33156 65560 33212
rect 65560 33156 65564 33212
rect 65500 33152 65564 33156
rect 64340 32668 64404 32672
rect 64340 32612 64344 32668
rect 64344 32612 64400 32668
rect 64400 32612 64404 32668
rect 64340 32608 64404 32612
rect 64420 32668 64484 32672
rect 64420 32612 64424 32668
rect 64424 32612 64480 32668
rect 64480 32612 64484 32668
rect 64420 32608 64484 32612
rect 64500 32668 64564 32672
rect 64500 32612 64504 32668
rect 64504 32612 64560 32668
rect 64560 32612 64564 32668
rect 64500 32608 64564 32612
rect 64580 32668 64644 32672
rect 64580 32612 64584 32668
rect 64584 32612 64640 32668
rect 64640 32612 64644 32668
rect 64580 32608 64644 32612
rect 65260 32124 65324 32128
rect 65260 32068 65264 32124
rect 65264 32068 65320 32124
rect 65320 32068 65324 32124
rect 65260 32064 65324 32068
rect 65340 32124 65404 32128
rect 65340 32068 65344 32124
rect 65344 32068 65400 32124
rect 65400 32068 65404 32124
rect 65340 32064 65404 32068
rect 65420 32124 65484 32128
rect 65420 32068 65424 32124
rect 65424 32068 65480 32124
rect 65480 32068 65484 32124
rect 65420 32064 65484 32068
rect 65500 32124 65564 32128
rect 65500 32068 65504 32124
rect 65504 32068 65560 32124
rect 65560 32068 65564 32124
rect 65500 32064 65564 32068
rect 64340 31580 64404 31584
rect 64340 31524 64344 31580
rect 64344 31524 64400 31580
rect 64400 31524 64404 31580
rect 64340 31520 64404 31524
rect 64420 31580 64484 31584
rect 64420 31524 64424 31580
rect 64424 31524 64480 31580
rect 64480 31524 64484 31580
rect 64420 31520 64484 31524
rect 64500 31580 64564 31584
rect 64500 31524 64504 31580
rect 64504 31524 64560 31580
rect 64560 31524 64564 31580
rect 64500 31520 64564 31524
rect 64580 31580 64644 31584
rect 64580 31524 64584 31580
rect 64584 31524 64640 31580
rect 64640 31524 64644 31580
rect 64580 31520 64644 31524
rect 65260 31036 65324 31040
rect 65260 30980 65264 31036
rect 65264 30980 65320 31036
rect 65320 30980 65324 31036
rect 65260 30976 65324 30980
rect 65340 31036 65404 31040
rect 65340 30980 65344 31036
rect 65344 30980 65400 31036
rect 65400 30980 65404 31036
rect 65340 30976 65404 30980
rect 65420 31036 65484 31040
rect 65420 30980 65424 31036
rect 65424 30980 65480 31036
rect 65480 30980 65484 31036
rect 65420 30976 65484 30980
rect 65500 31036 65564 31040
rect 65500 30980 65504 31036
rect 65504 30980 65560 31036
rect 65560 30980 65564 31036
rect 65500 30976 65564 30980
rect 64340 30492 64404 30496
rect 64340 30436 64344 30492
rect 64344 30436 64400 30492
rect 64400 30436 64404 30492
rect 64340 30432 64404 30436
rect 64420 30492 64484 30496
rect 64420 30436 64424 30492
rect 64424 30436 64480 30492
rect 64480 30436 64484 30492
rect 64420 30432 64484 30436
rect 64500 30492 64564 30496
rect 64500 30436 64504 30492
rect 64504 30436 64560 30492
rect 64560 30436 64564 30492
rect 64500 30432 64564 30436
rect 64580 30492 64644 30496
rect 64580 30436 64584 30492
rect 64584 30436 64640 30492
rect 64640 30436 64644 30492
rect 64580 30432 64644 30436
rect 65260 29948 65324 29952
rect 65260 29892 65264 29948
rect 65264 29892 65320 29948
rect 65320 29892 65324 29948
rect 65260 29888 65324 29892
rect 65340 29948 65404 29952
rect 65340 29892 65344 29948
rect 65344 29892 65400 29948
rect 65400 29892 65404 29948
rect 65340 29888 65404 29892
rect 65420 29948 65484 29952
rect 65420 29892 65424 29948
rect 65424 29892 65480 29948
rect 65480 29892 65484 29948
rect 65420 29888 65484 29892
rect 65500 29948 65564 29952
rect 65500 29892 65504 29948
rect 65504 29892 65560 29948
rect 65560 29892 65564 29948
rect 65500 29888 65564 29892
rect 64340 29404 64404 29408
rect 64340 29348 64344 29404
rect 64344 29348 64400 29404
rect 64400 29348 64404 29404
rect 64340 29344 64404 29348
rect 64420 29404 64484 29408
rect 64420 29348 64424 29404
rect 64424 29348 64480 29404
rect 64480 29348 64484 29404
rect 64420 29344 64484 29348
rect 64500 29404 64564 29408
rect 64500 29348 64504 29404
rect 64504 29348 64560 29404
rect 64560 29348 64564 29404
rect 64500 29344 64564 29348
rect 64580 29404 64644 29408
rect 64580 29348 64584 29404
rect 64584 29348 64640 29404
rect 64640 29348 64644 29404
rect 64580 29344 64644 29348
rect 62620 29178 62684 29242
rect 65260 28860 65324 28864
rect 65260 28804 65264 28860
rect 65264 28804 65320 28860
rect 65320 28804 65324 28860
rect 65260 28800 65324 28804
rect 65340 28860 65404 28864
rect 65340 28804 65344 28860
rect 65344 28804 65400 28860
rect 65400 28804 65404 28860
rect 65340 28800 65404 28804
rect 65420 28860 65484 28864
rect 65420 28804 65424 28860
rect 65424 28804 65480 28860
rect 65480 28804 65484 28860
rect 65420 28800 65484 28804
rect 65500 28860 65564 28864
rect 65500 28804 65504 28860
rect 65504 28804 65560 28860
rect 65560 28804 65564 28860
rect 65500 28800 65564 28804
rect 64340 28316 64404 28320
rect 64340 28260 64344 28316
rect 64344 28260 64400 28316
rect 64400 28260 64404 28316
rect 64340 28256 64404 28260
rect 64420 28316 64484 28320
rect 64420 28260 64424 28316
rect 64424 28260 64480 28316
rect 64480 28260 64484 28316
rect 64420 28256 64484 28260
rect 64500 28316 64564 28320
rect 64500 28260 64504 28316
rect 64504 28260 64560 28316
rect 64560 28260 64564 28316
rect 64500 28256 64564 28260
rect 64580 28316 64644 28320
rect 64580 28260 64584 28316
rect 64584 28260 64640 28316
rect 64640 28260 64644 28316
rect 64580 28256 64644 28260
rect 65260 27772 65324 27776
rect 65260 27716 65264 27772
rect 65264 27716 65320 27772
rect 65320 27716 65324 27772
rect 65260 27712 65324 27716
rect 65340 27772 65404 27776
rect 65340 27716 65344 27772
rect 65344 27716 65400 27772
rect 65400 27716 65404 27772
rect 65340 27712 65404 27716
rect 65420 27772 65484 27776
rect 65420 27716 65424 27772
rect 65424 27716 65480 27772
rect 65480 27716 65484 27772
rect 65420 27712 65484 27716
rect 65500 27772 65564 27776
rect 65500 27716 65504 27772
rect 65504 27716 65560 27772
rect 65560 27716 65564 27772
rect 65500 27712 65564 27716
rect 64340 27228 64404 27232
rect 64340 27172 64344 27228
rect 64344 27172 64400 27228
rect 64400 27172 64404 27228
rect 64340 27168 64404 27172
rect 64420 27228 64484 27232
rect 64420 27172 64424 27228
rect 64424 27172 64480 27228
rect 64480 27172 64484 27228
rect 64420 27168 64484 27172
rect 64500 27228 64564 27232
rect 64500 27172 64504 27228
rect 64504 27172 64560 27228
rect 64560 27172 64564 27228
rect 64500 27168 64564 27172
rect 64580 27228 64644 27232
rect 64580 27172 64584 27228
rect 64584 27172 64640 27228
rect 64640 27172 64644 27228
rect 64580 27168 64644 27172
rect 65260 26684 65324 26688
rect 65260 26628 65264 26684
rect 65264 26628 65320 26684
rect 65320 26628 65324 26684
rect 65260 26624 65324 26628
rect 65340 26684 65404 26688
rect 65340 26628 65344 26684
rect 65344 26628 65400 26684
rect 65400 26628 65404 26684
rect 65340 26624 65404 26628
rect 65420 26684 65484 26688
rect 65420 26628 65424 26684
rect 65424 26628 65480 26684
rect 65480 26628 65484 26684
rect 65420 26624 65484 26628
rect 65500 26684 65564 26688
rect 65500 26628 65504 26684
rect 65504 26628 65560 26684
rect 65560 26628 65564 26684
rect 65500 26624 65564 26628
rect 64340 26140 64404 26144
rect 64340 26084 64344 26140
rect 64344 26084 64400 26140
rect 64400 26084 64404 26140
rect 64340 26080 64404 26084
rect 64420 26140 64484 26144
rect 64420 26084 64424 26140
rect 64424 26084 64480 26140
rect 64480 26084 64484 26140
rect 64420 26080 64484 26084
rect 64500 26140 64564 26144
rect 64500 26084 64504 26140
rect 64504 26084 64560 26140
rect 64560 26084 64564 26140
rect 64500 26080 64564 26084
rect 64580 26140 64644 26144
rect 64580 26084 64584 26140
rect 64584 26084 64640 26140
rect 64640 26084 64644 26140
rect 64580 26080 64644 26084
rect 65260 25596 65324 25600
rect 65260 25540 65264 25596
rect 65264 25540 65320 25596
rect 65320 25540 65324 25596
rect 65260 25536 65324 25540
rect 65340 25596 65404 25600
rect 65340 25540 65344 25596
rect 65344 25540 65400 25596
rect 65400 25540 65404 25596
rect 65340 25536 65404 25540
rect 65420 25596 65484 25600
rect 65420 25540 65424 25596
rect 65424 25540 65480 25596
rect 65480 25540 65484 25596
rect 65420 25536 65484 25540
rect 65500 25596 65564 25600
rect 65500 25540 65504 25596
rect 65504 25540 65560 25596
rect 65560 25540 65564 25596
rect 65500 25536 65564 25540
rect 64340 25052 64404 25056
rect 64340 24996 64344 25052
rect 64344 24996 64400 25052
rect 64400 24996 64404 25052
rect 64340 24992 64404 24996
rect 64420 25052 64484 25056
rect 64420 24996 64424 25052
rect 64424 24996 64480 25052
rect 64480 24996 64484 25052
rect 64420 24992 64484 24996
rect 64500 25052 64564 25056
rect 64500 24996 64504 25052
rect 64504 24996 64560 25052
rect 64560 24996 64564 25052
rect 64500 24992 64564 24996
rect 64580 25052 64644 25056
rect 64580 24996 64584 25052
rect 64584 24996 64640 25052
rect 64640 24996 64644 25052
rect 64580 24992 64644 24996
rect 65260 24508 65324 24512
rect 65260 24452 65264 24508
rect 65264 24452 65320 24508
rect 65320 24452 65324 24508
rect 65260 24448 65324 24452
rect 65340 24508 65404 24512
rect 65340 24452 65344 24508
rect 65344 24452 65400 24508
rect 65400 24452 65404 24508
rect 65340 24448 65404 24452
rect 65420 24508 65484 24512
rect 65420 24452 65424 24508
rect 65424 24452 65480 24508
rect 65480 24452 65484 24508
rect 65420 24448 65484 24452
rect 65500 24508 65564 24512
rect 65500 24452 65504 24508
rect 65504 24452 65560 24508
rect 65560 24452 65564 24508
rect 65500 24448 65564 24452
rect 64340 23964 64404 23968
rect 64340 23908 64344 23964
rect 64344 23908 64400 23964
rect 64400 23908 64404 23964
rect 64340 23904 64404 23908
rect 64420 23964 64484 23968
rect 64420 23908 64424 23964
rect 64424 23908 64480 23964
rect 64480 23908 64484 23964
rect 64420 23904 64484 23908
rect 64500 23964 64564 23968
rect 64500 23908 64504 23964
rect 64504 23908 64560 23964
rect 64560 23908 64564 23964
rect 64500 23904 64564 23908
rect 64580 23964 64644 23968
rect 64580 23908 64584 23964
rect 64584 23908 64640 23964
rect 64640 23908 64644 23964
rect 64580 23904 64644 23908
rect 65260 23420 65324 23424
rect 65260 23364 65264 23420
rect 65264 23364 65320 23420
rect 65320 23364 65324 23420
rect 65260 23360 65324 23364
rect 65340 23420 65404 23424
rect 65340 23364 65344 23420
rect 65344 23364 65400 23420
rect 65400 23364 65404 23420
rect 65340 23360 65404 23364
rect 65420 23420 65484 23424
rect 65420 23364 65424 23420
rect 65424 23364 65480 23420
rect 65480 23364 65484 23420
rect 65420 23360 65484 23364
rect 65500 23420 65564 23424
rect 65500 23364 65504 23420
rect 65504 23364 65560 23420
rect 65560 23364 65564 23420
rect 65500 23360 65564 23364
rect 64340 22876 64404 22880
rect 64340 22820 64344 22876
rect 64344 22820 64400 22876
rect 64400 22820 64404 22876
rect 64340 22816 64404 22820
rect 64420 22876 64484 22880
rect 64420 22820 64424 22876
rect 64424 22820 64480 22876
rect 64480 22820 64484 22876
rect 64420 22816 64484 22820
rect 64500 22876 64564 22880
rect 64500 22820 64504 22876
rect 64504 22820 64560 22876
rect 64560 22820 64564 22876
rect 64500 22816 64564 22820
rect 64580 22876 64644 22880
rect 64580 22820 64584 22876
rect 64584 22820 64640 22876
rect 64640 22820 64644 22876
rect 64580 22816 64644 22820
rect 65260 22332 65324 22336
rect 65260 22276 65264 22332
rect 65264 22276 65320 22332
rect 65320 22276 65324 22332
rect 65260 22272 65324 22276
rect 65340 22332 65404 22336
rect 65340 22276 65344 22332
rect 65344 22276 65400 22332
rect 65400 22276 65404 22332
rect 65340 22272 65404 22276
rect 65420 22332 65484 22336
rect 65420 22276 65424 22332
rect 65424 22276 65480 22332
rect 65480 22276 65484 22332
rect 65420 22272 65484 22276
rect 65500 22332 65564 22336
rect 65500 22276 65504 22332
rect 65504 22276 65560 22332
rect 65560 22276 65564 22332
rect 65500 22272 65564 22276
rect 64340 21788 64404 21792
rect 64340 21732 64344 21788
rect 64344 21732 64400 21788
rect 64400 21732 64404 21788
rect 64340 21728 64404 21732
rect 64420 21788 64484 21792
rect 64420 21732 64424 21788
rect 64424 21732 64480 21788
rect 64480 21732 64484 21788
rect 64420 21728 64484 21732
rect 64500 21788 64564 21792
rect 64500 21732 64504 21788
rect 64504 21732 64560 21788
rect 64560 21732 64564 21788
rect 64500 21728 64564 21732
rect 64580 21788 64644 21792
rect 64580 21732 64584 21788
rect 64584 21732 64640 21788
rect 64640 21732 64644 21788
rect 64580 21728 64644 21732
rect 65260 21244 65324 21248
rect 65260 21188 65264 21244
rect 65264 21188 65320 21244
rect 65320 21188 65324 21244
rect 65260 21184 65324 21188
rect 65340 21244 65404 21248
rect 65340 21188 65344 21244
rect 65344 21188 65400 21244
rect 65400 21188 65404 21244
rect 65340 21184 65404 21188
rect 65420 21244 65484 21248
rect 65420 21188 65424 21244
rect 65424 21188 65480 21244
rect 65480 21188 65484 21244
rect 65420 21184 65484 21188
rect 65500 21244 65564 21248
rect 65500 21188 65504 21244
rect 65504 21188 65560 21244
rect 65560 21188 65564 21244
rect 65500 21184 65564 21188
rect 64340 20700 64404 20704
rect 64340 20644 64344 20700
rect 64344 20644 64400 20700
rect 64400 20644 64404 20700
rect 64340 20640 64404 20644
rect 64420 20700 64484 20704
rect 64420 20644 64424 20700
rect 64424 20644 64480 20700
rect 64480 20644 64484 20700
rect 64420 20640 64484 20644
rect 64500 20700 64564 20704
rect 64500 20644 64504 20700
rect 64504 20644 64560 20700
rect 64560 20644 64564 20700
rect 64500 20640 64564 20644
rect 64580 20700 64644 20704
rect 64580 20644 64584 20700
rect 64584 20644 64640 20700
rect 64640 20644 64644 20700
rect 64580 20640 64644 20644
rect 65260 20156 65324 20160
rect 65260 20100 65264 20156
rect 65264 20100 65320 20156
rect 65320 20100 65324 20156
rect 65260 20096 65324 20100
rect 65340 20156 65404 20160
rect 65340 20100 65344 20156
rect 65344 20100 65400 20156
rect 65400 20100 65404 20156
rect 65340 20096 65404 20100
rect 65420 20156 65484 20160
rect 65420 20100 65424 20156
rect 65424 20100 65480 20156
rect 65480 20100 65484 20156
rect 65420 20096 65484 20100
rect 65500 20156 65564 20160
rect 65500 20100 65504 20156
rect 65504 20100 65560 20156
rect 65560 20100 65564 20156
rect 65500 20096 65564 20100
rect 64340 19612 64404 19616
rect 64340 19556 64344 19612
rect 64344 19556 64400 19612
rect 64400 19556 64404 19612
rect 64340 19552 64404 19556
rect 64420 19612 64484 19616
rect 64420 19556 64424 19612
rect 64424 19556 64480 19612
rect 64480 19556 64484 19612
rect 64420 19552 64484 19556
rect 64500 19612 64564 19616
rect 64500 19556 64504 19612
rect 64504 19556 64560 19612
rect 64560 19556 64564 19612
rect 64500 19552 64564 19556
rect 64580 19612 64644 19616
rect 64580 19556 64584 19612
rect 64584 19556 64640 19612
rect 64640 19556 64644 19612
rect 64580 19552 64644 19556
rect 65260 19068 65324 19072
rect 65260 19012 65264 19068
rect 65264 19012 65320 19068
rect 65320 19012 65324 19068
rect 65260 19008 65324 19012
rect 65340 19068 65404 19072
rect 65340 19012 65344 19068
rect 65344 19012 65400 19068
rect 65400 19012 65404 19068
rect 65340 19008 65404 19012
rect 65420 19068 65484 19072
rect 65420 19012 65424 19068
rect 65424 19012 65480 19068
rect 65480 19012 65484 19068
rect 65420 19008 65484 19012
rect 65500 19068 65564 19072
rect 65500 19012 65504 19068
rect 65504 19012 65560 19068
rect 65560 19012 65564 19068
rect 65500 19008 65564 19012
rect 64340 18524 64404 18528
rect 64340 18468 64344 18524
rect 64344 18468 64400 18524
rect 64400 18468 64404 18524
rect 64340 18464 64404 18468
rect 64420 18524 64484 18528
rect 64420 18468 64424 18524
rect 64424 18468 64480 18524
rect 64480 18468 64484 18524
rect 64420 18464 64484 18468
rect 64500 18524 64564 18528
rect 64500 18468 64504 18524
rect 64504 18468 64560 18524
rect 64560 18468 64564 18524
rect 64500 18464 64564 18468
rect 64580 18524 64644 18528
rect 64580 18468 64584 18524
rect 64584 18468 64640 18524
rect 64640 18468 64644 18524
rect 64580 18464 64644 18468
rect 65260 17980 65324 17984
rect 65260 17924 65264 17980
rect 65264 17924 65320 17980
rect 65320 17924 65324 17980
rect 65260 17920 65324 17924
rect 65340 17980 65404 17984
rect 65340 17924 65344 17980
rect 65344 17924 65400 17980
rect 65400 17924 65404 17980
rect 65340 17920 65404 17924
rect 65420 17980 65484 17984
rect 65420 17924 65424 17980
rect 65424 17924 65480 17980
rect 65480 17924 65484 17980
rect 65420 17920 65484 17924
rect 65500 17980 65564 17984
rect 65500 17924 65504 17980
rect 65504 17924 65560 17980
rect 65560 17924 65564 17980
rect 65500 17920 65564 17924
rect 64340 17436 64404 17440
rect 64340 17380 64344 17436
rect 64344 17380 64400 17436
rect 64400 17380 64404 17436
rect 64340 17376 64404 17380
rect 64420 17436 64484 17440
rect 64420 17380 64424 17436
rect 64424 17380 64480 17436
rect 64480 17380 64484 17436
rect 64420 17376 64484 17380
rect 64500 17436 64564 17440
rect 64500 17380 64504 17436
rect 64504 17380 64560 17436
rect 64560 17380 64564 17436
rect 64500 17376 64564 17380
rect 64580 17436 64644 17440
rect 64580 17380 64584 17436
rect 64584 17380 64640 17436
rect 64640 17380 64644 17436
rect 64580 17376 64644 17380
rect 65260 16892 65324 16896
rect 65260 16836 65264 16892
rect 65264 16836 65320 16892
rect 65320 16836 65324 16892
rect 65260 16832 65324 16836
rect 65340 16892 65404 16896
rect 65340 16836 65344 16892
rect 65344 16836 65400 16892
rect 65400 16836 65404 16892
rect 65340 16832 65404 16836
rect 65420 16892 65484 16896
rect 65420 16836 65424 16892
rect 65424 16836 65480 16892
rect 65480 16836 65484 16892
rect 65420 16832 65484 16836
rect 65500 16892 65564 16896
rect 65500 16836 65504 16892
rect 65504 16836 65560 16892
rect 65560 16836 65564 16892
rect 65500 16832 65564 16836
rect 64340 16348 64404 16352
rect 64340 16292 64344 16348
rect 64344 16292 64400 16348
rect 64400 16292 64404 16348
rect 64340 16288 64404 16292
rect 64420 16348 64484 16352
rect 64420 16292 64424 16348
rect 64424 16292 64480 16348
rect 64480 16292 64484 16348
rect 64420 16288 64484 16292
rect 64500 16348 64564 16352
rect 64500 16292 64504 16348
rect 64504 16292 64560 16348
rect 64560 16292 64564 16348
rect 64500 16288 64564 16292
rect 64580 16348 64644 16352
rect 64580 16292 64584 16348
rect 64584 16292 64640 16348
rect 64640 16292 64644 16348
rect 64580 16288 64644 16292
rect 65260 15804 65324 15808
rect 65260 15748 65264 15804
rect 65264 15748 65320 15804
rect 65320 15748 65324 15804
rect 65260 15744 65324 15748
rect 65340 15804 65404 15808
rect 65340 15748 65344 15804
rect 65344 15748 65400 15804
rect 65400 15748 65404 15804
rect 65340 15744 65404 15748
rect 65420 15804 65484 15808
rect 65420 15748 65424 15804
rect 65424 15748 65480 15804
rect 65480 15748 65484 15804
rect 65420 15744 65484 15748
rect 65500 15804 65564 15808
rect 65500 15748 65504 15804
rect 65504 15748 65560 15804
rect 65560 15748 65564 15804
rect 65500 15744 65564 15748
rect 63356 15268 63420 15332
rect 64340 15260 64404 15264
rect 64340 15204 64344 15260
rect 64344 15204 64400 15260
rect 64400 15204 64404 15260
rect 64340 15200 64404 15204
rect 64420 15260 64484 15264
rect 64420 15204 64424 15260
rect 64424 15204 64480 15260
rect 64480 15204 64484 15260
rect 64420 15200 64484 15204
rect 64500 15260 64564 15264
rect 64500 15204 64504 15260
rect 64504 15204 64560 15260
rect 64560 15204 64564 15260
rect 64500 15200 64564 15204
rect 64580 15260 64644 15264
rect 64580 15204 64584 15260
rect 64584 15204 64640 15260
rect 64640 15204 64644 15260
rect 64580 15200 64644 15204
rect 65260 14716 65324 14720
rect 65260 14660 65264 14716
rect 65264 14660 65320 14716
rect 65320 14660 65324 14716
rect 65260 14656 65324 14660
rect 65340 14716 65404 14720
rect 65340 14660 65344 14716
rect 65344 14660 65400 14716
rect 65400 14660 65404 14716
rect 65340 14656 65404 14660
rect 65420 14716 65484 14720
rect 65420 14660 65424 14716
rect 65424 14660 65480 14716
rect 65480 14660 65484 14716
rect 65420 14656 65484 14660
rect 65500 14716 65564 14720
rect 65500 14660 65504 14716
rect 65504 14660 65560 14716
rect 65560 14660 65564 14716
rect 65500 14656 65564 14660
rect 64340 14172 64404 14176
rect 64340 14116 64344 14172
rect 64344 14116 64400 14172
rect 64400 14116 64404 14172
rect 64340 14112 64404 14116
rect 64420 14172 64484 14176
rect 64420 14116 64424 14172
rect 64424 14116 64480 14172
rect 64480 14116 64484 14172
rect 64420 14112 64484 14116
rect 64500 14172 64564 14176
rect 64500 14116 64504 14172
rect 64504 14116 64560 14172
rect 64560 14116 64564 14172
rect 64500 14112 64564 14116
rect 64580 14172 64644 14176
rect 64580 14116 64584 14172
rect 64584 14116 64640 14172
rect 64640 14116 64644 14172
rect 64580 14112 64644 14116
rect 65260 13628 65324 13632
rect 65260 13572 65264 13628
rect 65264 13572 65320 13628
rect 65320 13572 65324 13628
rect 65260 13568 65324 13572
rect 65340 13628 65404 13632
rect 65340 13572 65344 13628
rect 65344 13572 65400 13628
rect 65400 13572 65404 13628
rect 65340 13568 65404 13572
rect 65420 13628 65484 13632
rect 65420 13572 65424 13628
rect 65424 13572 65480 13628
rect 65480 13572 65484 13628
rect 65420 13568 65484 13572
rect 65500 13628 65564 13632
rect 65500 13572 65504 13628
rect 65504 13572 65560 13628
rect 65560 13572 65564 13628
rect 65500 13568 65564 13572
rect 64340 13084 64404 13088
rect 64340 13028 64344 13084
rect 64344 13028 64400 13084
rect 64400 13028 64404 13084
rect 64340 13024 64404 13028
rect 64420 13084 64484 13088
rect 64420 13028 64424 13084
rect 64424 13028 64480 13084
rect 64480 13028 64484 13084
rect 64420 13024 64484 13028
rect 64500 13084 64564 13088
rect 64500 13028 64504 13084
rect 64504 13028 64560 13084
rect 64560 13028 64564 13084
rect 64500 13024 64564 13028
rect 64580 13084 64644 13088
rect 64580 13028 64584 13084
rect 64584 13028 64640 13084
rect 64640 13028 64644 13084
rect 64580 13024 64644 13028
rect 65260 12540 65324 12544
rect 65260 12484 65264 12540
rect 65264 12484 65320 12540
rect 65320 12484 65324 12540
rect 65260 12480 65324 12484
rect 65340 12540 65404 12544
rect 65340 12484 65344 12540
rect 65344 12484 65400 12540
rect 65400 12484 65404 12540
rect 65340 12480 65404 12484
rect 65420 12540 65484 12544
rect 65420 12484 65424 12540
rect 65424 12484 65480 12540
rect 65480 12484 65484 12540
rect 65420 12480 65484 12484
rect 65500 12540 65564 12544
rect 65500 12484 65504 12540
rect 65504 12484 65560 12540
rect 65560 12484 65564 12540
rect 65500 12480 65564 12484
rect 64340 11996 64404 12000
rect 64340 11940 64344 11996
rect 64344 11940 64400 11996
rect 64400 11940 64404 11996
rect 64340 11936 64404 11940
rect 64420 11996 64484 12000
rect 64420 11940 64424 11996
rect 64424 11940 64480 11996
rect 64480 11940 64484 11996
rect 64420 11936 64484 11940
rect 64500 11996 64564 12000
rect 64500 11940 64504 11996
rect 64504 11940 64560 11996
rect 64560 11940 64564 11996
rect 64500 11936 64564 11940
rect 64580 11996 64644 12000
rect 64580 11940 64584 11996
rect 64584 11940 64640 11996
rect 64640 11940 64644 11996
rect 64580 11936 64644 11940
rect 65260 11452 65324 11456
rect 65260 11396 65264 11452
rect 65264 11396 65320 11452
rect 65320 11396 65324 11452
rect 65260 11392 65324 11396
rect 65340 11452 65404 11456
rect 65340 11396 65344 11452
rect 65344 11396 65400 11452
rect 65400 11396 65404 11452
rect 65340 11392 65404 11396
rect 65420 11452 65484 11456
rect 65420 11396 65424 11452
rect 65424 11396 65480 11452
rect 65480 11396 65484 11452
rect 65420 11392 65484 11396
rect 65500 11452 65564 11456
rect 65500 11396 65504 11452
rect 65504 11396 65560 11452
rect 65560 11396 65564 11452
rect 65500 11392 65564 11396
rect 64340 10908 64404 10912
rect 64340 10852 64344 10908
rect 64344 10852 64400 10908
rect 64400 10852 64404 10908
rect 64340 10848 64404 10852
rect 64420 10908 64484 10912
rect 64420 10852 64424 10908
rect 64424 10852 64480 10908
rect 64480 10852 64484 10908
rect 64420 10848 64484 10852
rect 64500 10908 64564 10912
rect 64500 10852 64504 10908
rect 64504 10852 64560 10908
rect 64560 10852 64564 10908
rect 64500 10848 64564 10852
rect 64580 10908 64644 10912
rect 64580 10852 64584 10908
rect 64584 10852 64640 10908
rect 64640 10852 64644 10908
rect 64580 10848 64644 10852
rect 65260 10364 65324 10368
rect 65260 10308 65264 10364
rect 65264 10308 65320 10364
rect 65320 10308 65324 10364
rect 65260 10304 65324 10308
rect 65340 10364 65404 10368
rect 65340 10308 65344 10364
rect 65344 10308 65400 10364
rect 65400 10308 65404 10364
rect 65340 10304 65404 10308
rect 65420 10364 65484 10368
rect 65420 10308 65424 10364
rect 65424 10308 65480 10364
rect 65480 10308 65484 10364
rect 65420 10304 65484 10308
rect 65500 10364 65564 10368
rect 65500 10308 65504 10364
rect 65504 10308 65560 10364
rect 65560 10308 65564 10364
rect 65500 10304 65564 10308
rect 64340 9820 64404 9824
rect 64340 9764 64344 9820
rect 64344 9764 64400 9820
rect 64400 9764 64404 9820
rect 64340 9760 64404 9764
rect 64420 9820 64484 9824
rect 64420 9764 64424 9820
rect 64424 9764 64480 9820
rect 64480 9764 64484 9820
rect 64420 9760 64484 9764
rect 64500 9820 64564 9824
rect 64500 9764 64504 9820
rect 64504 9764 64560 9820
rect 64560 9764 64564 9820
rect 64500 9760 64564 9764
rect 64580 9820 64644 9824
rect 64580 9764 64584 9820
rect 64584 9764 64640 9820
rect 64640 9764 64644 9820
rect 64580 9760 64644 9764
rect 65260 9276 65324 9280
rect 65260 9220 65264 9276
rect 65264 9220 65320 9276
rect 65320 9220 65324 9276
rect 65260 9216 65324 9220
rect 65340 9276 65404 9280
rect 65340 9220 65344 9276
rect 65344 9220 65400 9276
rect 65400 9220 65404 9276
rect 65340 9216 65404 9220
rect 65420 9276 65484 9280
rect 65420 9220 65424 9276
rect 65424 9220 65480 9276
rect 65480 9220 65484 9276
rect 65420 9216 65484 9220
rect 65500 9276 65564 9280
rect 65500 9220 65504 9276
rect 65504 9220 65560 9276
rect 65560 9220 65564 9276
rect 65500 9216 65564 9220
rect 64340 8732 64404 8736
rect 64340 8676 64344 8732
rect 64344 8676 64400 8732
rect 64400 8676 64404 8732
rect 64340 8672 64404 8676
rect 64420 8732 64484 8736
rect 64420 8676 64424 8732
rect 64424 8676 64480 8732
rect 64480 8676 64484 8732
rect 64420 8672 64484 8676
rect 64500 8732 64564 8736
rect 64500 8676 64504 8732
rect 64504 8676 64560 8732
rect 64560 8676 64564 8732
rect 64500 8672 64564 8676
rect 64580 8732 64644 8736
rect 64580 8676 64584 8732
rect 64584 8676 64640 8732
rect 64640 8676 64644 8732
rect 64580 8672 64644 8676
rect 65260 8188 65324 8192
rect 65260 8132 65264 8188
rect 65264 8132 65320 8188
rect 65320 8132 65324 8188
rect 65260 8128 65324 8132
rect 65340 8188 65404 8192
rect 65340 8132 65344 8188
rect 65344 8132 65400 8188
rect 65400 8132 65404 8188
rect 65340 8128 65404 8132
rect 65420 8188 65484 8192
rect 65420 8132 65424 8188
rect 65424 8132 65480 8188
rect 65480 8132 65484 8188
rect 65420 8128 65484 8132
rect 65500 8188 65564 8192
rect 65500 8132 65504 8188
rect 65504 8132 65560 8188
rect 65560 8132 65564 8188
rect 65500 8128 65564 8132
rect 64340 7644 64404 7648
rect 64340 7588 64344 7644
rect 64344 7588 64400 7644
rect 64400 7588 64404 7644
rect 64340 7584 64404 7588
rect 64420 7644 64484 7648
rect 64420 7588 64424 7644
rect 64424 7588 64480 7644
rect 64480 7588 64484 7644
rect 64420 7584 64484 7588
rect 64500 7644 64564 7648
rect 64500 7588 64504 7644
rect 64504 7588 64560 7644
rect 64560 7588 64564 7644
rect 64500 7584 64564 7588
rect 64580 7644 64644 7648
rect 64580 7588 64584 7644
rect 64584 7588 64640 7644
rect 64640 7588 64644 7644
rect 64580 7584 64644 7588
rect 65260 7100 65324 7104
rect 65260 7044 65264 7100
rect 65264 7044 65320 7100
rect 65320 7044 65324 7100
rect 65260 7040 65324 7044
rect 65340 7100 65404 7104
rect 65340 7044 65344 7100
rect 65344 7044 65400 7100
rect 65400 7044 65404 7100
rect 65340 7040 65404 7044
rect 65420 7100 65484 7104
rect 65420 7044 65424 7100
rect 65424 7044 65480 7100
rect 65480 7044 65484 7100
rect 65420 7040 65484 7044
rect 65500 7100 65564 7104
rect 65500 7044 65504 7100
rect 65504 7044 65560 7100
rect 65560 7044 65564 7100
rect 65500 7040 65564 7044
rect 64340 6556 64404 6560
rect 64340 6500 64344 6556
rect 64344 6500 64400 6556
rect 64400 6500 64404 6556
rect 64340 6496 64404 6500
rect 64420 6556 64484 6560
rect 64420 6500 64424 6556
rect 64424 6500 64480 6556
rect 64480 6500 64484 6556
rect 64420 6496 64484 6500
rect 64500 6556 64564 6560
rect 64500 6500 64504 6556
rect 64504 6500 64560 6556
rect 64560 6500 64564 6556
rect 64500 6496 64564 6500
rect 64580 6556 64644 6560
rect 64580 6500 64584 6556
rect 64584 6500 64640 6556
rect 64640 6500 64644 6556
rect 64580 6496 64644 6500
rect 63908 6020 63972 6084
rect 65260 6012 65324 6016
rect 65260 5956 65264 6012
rect 65264 5956 65320 6012
rect 65320 5956 65324 6012
rect 65260 5952 65324 5956
rect 65340 6012 65404 6016
rect 65340 5956 65344 6012
rect 65344 5956 65400 6012
rect 65400 5956 65404 6012
rect 65340 5952 65404 5956
rect 65420 6012 65484 6016
rect 65420 5956 65424 6012
rect 65424 5956 65480 6012
rect 65480 5956 65484 6012
rect 65420 5952 65484 5956
rect 65500 6012 65564 6016
rect 65500 5956 65504 6012
rect 65504 5956 65560 6012
rect 65560 5956 65564 6012
rect 65500 5952 65564 5956
rect 64092 5944 64156 5948
rect 64092 5888 64142 5944
rect 64142 5888 64156 5944
rect 64092 5884 64156 5888
rect 64340 5468 64404 5472
rect 64340 5412 64344 5468
rect 64344 5412 64400 5468
rect 64400 5412 64404 5468
rect 64340 5408 64404 5412
rect 64420 5468 64484 5472
rect 64420 5412 64424 5468
rect 64424 5412 64480 5468
rect 64480 5412 64484 5468
rect 64420 5408 64484 5412
rect 64500 5468 64564 5472
rect 64500 5412 64504 5468
rect 64504 5412 64560 5468
rect 64560 5412 64564 5468
rect 64500 5408 64564 5412
rect 64580 5468 64644 5472
rect 64580 5412 64584 5468
rect 64584 5412 64640 5468
rect 64640 5412 64644 5468
rect 64580 5408 64644 5412
rect 65260 4924 65324 4928
rect 65260 4868 65264 4924
rect 65264 4868 65320 4924
rect 65320 4868 65324 4924
rect 65260 4864 65324 4868
rect 65340 4924 65404 4928
rect 65340 4868 65344 4924
rect 65344 4868 65400 4924
rect 65400 4868 65404 4924
rect 65340 4864 65404 4868
rect 65420 4924 65484 4928
rect 65420 4868 65424 4924
rect 65424 4868 65480 4924
rect 65480 4868 65484 4924
rect 65420 4864 65484 4868
rect 65500 4924 65564 4928
rect 65500 4868 65504 4924
rect 65504 4868 65560 4924
rect 65560 4868 65564 4924
rect 65500 4864 65564 4868
rect 64340 4380 64404 4384
rect 64340 4324 64344 4380
rect 64344 4324 64400 4380
rect 64400 4324 64404 4380
rect 64340 4320 64404 4324
rect 64420 4380 64484 4384
rect 64420 4324 64424 4380
rect 64424 4324 64480 4380
rect 64480 4324 64484 4380
rect 64420 4320 64484 4324
rect 64500 4380 64564 4384
rect 64500 4324 64504 4380
rect 64504 4324 64560 4380
rect 64560 4324 64564 4380
rect 64500 4320 64564 4324
rect 64580 4380 64644 4384
rect 64580 4324 64584 4380
rect 64584 4324 64640 4380
rect 64640 4324 64644 4380
rect 64580 4320 64644 4324
rect 65260 3836 65324 3840
rect 65260 3780 65264 3836
rect 65264 3780 65320 3836
rect 65320 3780 65324 3836
rect 65260 3776 65324 3780
rect 65340 3836 65404 3840
rect 65340 3780 65344 3836
rect 65344 3780 65400 3836
rect 65400 3780 65404 3836
rect 65340 3776 65404 3780
rect 65420 3836 65484 3840
rect 65420 3780 65424 3836
rect 65424 3780 65480 3836
rect 65480 3780 65484 3836
rect 65420 3776 65484 3780
rect 65500 3836 65564 3840
rect 65500 3780 65504 3836
rect 65504 3780 65560 3836
rect 65560 3780 65564 3836
rect 65500 3776 65564 3780
rect 64340 3292 64404 3296
rect 64340 3236 64344 3292
rect 64344 3236 64400 3292
rect 64400 3236 64404 3292
rect 64340 3232 64404 3236
rect 64420 3292 64484 3296
rect 64420 3236 64424 3292
rect 64424 3236 64480 3292
rect 64480 3236 64484 3292
rect 64420 3232 64484 3236
rect 64500 3292 64564 3296
rect 64500 3236 64504 3292
rect 64504 3236 64560 3292
rect 64560 3236 64564 3292
rect 64500 3232 64564 3236
rect 64580 3292 64644 3296
rect 64580 3236 64584 3292
rect 64584 3236 64640 3292
rect 64640 3236 64644 3292
rect 64580 3232 64644 3236
rect 65260 2748 65324 2752
rect 65260 2692 65264 2748
rect 65264 2692 65320 2748
rect 65320 2692 65324 2748
rect 65260 2688 65324 2692
rect 65340 2748 65404 2752
rect 65340 2692 65344 2748
rect 65344 2692 65400 2748
rect 65400 2692 65404 2748
rect 65340 2688 65404 2692
rect 65420 2748 65484 2752
rect 65420 2692 65424 2748
rect 65424 2692 65480 2748
rect 65480 2692 65484 2748
rect 65420 2688 65484 2692
rect 65500 2748 65564 2752
rect 65500 2692 65504 2748
rect 65504 2692 65560 2748
rect 65560 2692 65564 2748
rect 65500 2688 65564 2692
rect 64340 2204 64404 2208
rect 64340 2148 64344 2204
rect 64344 2148 64400 2204
rect 64400 2148 64404 2204
rect 64340 2144 64404 2148
rect 64420 2204 64484 2208
rect 64420 2148 64424 2204
rect 64424 2148 64480 2204
rect 64480 2148 64484 2204
rect 64420 2144 64484 2148
rect 64500 2204 64564 2208
rect 64500 2148 64504 2204
rect 64504 2148 64560 2204
rect 64560 2148 64564 2204
rect 64500 2144 64564 2148
rect 64580 2204 64644 2208
rect 64580 2148 64584 2204
rect 64584 2148 64640 2204
rect 64640 2148 64644 2204
rect 64580 2144 64644 2148
rect 63724 1940 63788 2004
rect 48941 1864 49005 1868
rect 48941 1808 48962 1864
rect 48962 1808 49005 1864
rect 48941 1804 49005 1808
rect 49217 1864 49281 1868
rect 49217 1808 49238 1864
rect 49238 1808 49281 1864
rect 49217 1804 49281 1808
rect 49674 1864 49738 1868
rect 49674 1808 49698 1864
rect 49698 1808 49738 1864
rect 49674 1804 49738 1808
rect 49372 1668 49436 1732
rect 65260 1660 65324 1664
rect 65260 1604 65264 1660
rect 65264 1604 65320 1660
rect 65320 1604 65324 1660
rect 65260 1600 65324 1604
rect 65340 1660 65404 1664
rect 65340 1604 65344 1660
rect 65344 1604 65400 1660
rect 65400 1604 65404 1660
rect 65340 1600 65404 1604
rect 65420 1660 65484 1664
rect 65420 1604 65424 1660
rect 65424 1604 65480 1660
rect 65480 1604 65484 1660
rect 65420 1600 65484 1604
rect 65500 1660 65564 1664
rect 65500 1604 65504 1660
rect 65504 1604 65560 1660
rect 65560 1604 65564 1660
rect 65500 1600 65564 1604
rect 49079 1532 49143 1596
rect 49924 1260 49988 1324
rect 64340 1116 64404 1120
rect 64340 1060 64344 1116
rect 64344 1060 64400 1116
rect 64400 1060 64404 1116
rect 64340 1056 64404 1060
rect 64420 1116 64484 1120
rect 64420 1060 64424 1116
rect 64424 1060 64480 1116
rect 64480 1060 64484 1116
rect 64420 1056 64484 1060
rect 64500 1116 64564 1120
rect 64500 1060 64504 1116
rect 64504 1060 64560 1116
rect 64560 1060 64564 1116
rect 64500 1056 64564 1060
rect 64580 1116 64644 1120
rect 64580 1060 64584 1116
rect 64584 1060 64640 1116
rect 64640 1060 64644 1116
rect 64580 1056 64644 1060
rect 65260 572 65324 576
rect 65260 516 65264 572
rect 65264 516 65320 572
rect 65320 516 65324 572
rect 65260 512 65324 516
rect 65340 572 65404 576
rect 65340 516 65344 572
rect 65344 516 65400 572
rect 65400 516 65404 572
rect 65340 512 65404 516
rect 65420 572 65484 576
rect 65420 516 65424 572
rect 65424 516 65480 572
rect 65480 516 65484 572
rect 65420 512 65484 516
rect 65500 572 65564 576
rect 65500 516 65504 572
rect 65504 516 65560 572
rect 65560 516 65564 572
rect 65500 512 65564 516
<< metal4 >>
rect 1992 44640 2312 44656
rect 1992 44576 2000 44640
rect 2064 44576 2080 44640
rect 2144 44576 2160 44640
rect 2224 44576 2240 44640
rect 2304 44576 2312 44640
rect 1992 43552 2312 44576
rect 1992 43488 2000 43552
rect 2064 43488 2080 43552
rect 2144 43488 2160 43552
rect 2224 43488 2240 43552
rect 2304 43488 2312 43552
rect 1992 42464 2312 43488
rect 1992 42400 2000 42464
rect 2064 42400 2080 42464
rect 2144 42400 2160 42464
rect 2224 42400 2240 42464
rect 2304 42400 2312 42464
rect 1992 41376 2312 42400
rect 1992 41312 2000 41376
rect 2064 41312 2080 41376
rect 2144 41312 2160 41376
rect 2224 41312 2240 41376
rect 2304 41312 2312 41376
rect 1992 40288 2312 41312
rect 1992 40224 2000 40288
rect 2064 40224 2080 40288
rect 2144 40224 2160 40288
rect 2224 40224 2240 40288
rect 2304 40224 2312 40288
rect 1992 39200 2312 40224
rect 1992 39136 2000 39200
rect 2064 39136 2080 39200
rect 2144 39136 2160 39200
rect 2224 39136 2240 39200
rect 2304 39136 2312 39200
rect 1992 38112 2312 39136
rect 1992 38048 2000 38112
rect 2064 38048 2080 38112
rect 2144 38048 2160 38112
rect 2224 38048 2240 38112
rect 2304 38048 2312 38112
rect 1992 37024 2312 38048
rect 1992 36960 2000 37024
rect 2064 36960 2080 37024
rect 2144 36960 2160 37024
rect 2224 36960 2240 37024
rect 2304 36960 2312 37024
rect 1992 35492 2312 36960
rect 1992 35428 2000 35492
rect 2064 35428 2080 35492
rect 2144 35428 2160 35492
rect 2224 35428 2240 35492
rect 2304 35428 2312 35492
rect 1992 35412 2312 35428
rect 1992 35348 2000 35412
rect 2064 35348 2080 35412
rect 2144 35348 2160 35412
rect 2224 35348 2240 35412
rect 2304 35348 2312 35412
rect 1992 35332 2312 35348
rect 1992 35268 2000 35332
rect 2064 35268 2080 35332
rect 2144 35268 2160 35332
rect 2224 35268 2240 35332
rect 2304 35268 2312 35332
rect 1992 35252 2312 35268
rect 1992 35188 2000 35252
rect 2064 35188 2080 35252
rect 2144 35188 2160 35252
rect 2224 35188 2240 35252
rect 2304 35188 2312 35252
rect 1992 34208 2312 35188
rect 2912 44096 3232 44656
rect 6134 44573 6194 45152
rect 6686 44573 6746 45152
rect 7238 44573 7298 45152
rect 7790 44573 7850 45152
rect 8342 44573 8402 45152
rect 8894 44573 8954 45152
rect 9446 44573 9506 45152
rect 9998 44573 10058 45152
rect 10550 44573 10610 45152
rect 6131 44572 6197 44573
rect 6131 44508 6132 44572
rect 6196 44508 6197 44572
rect 6131 44507 6197 44508
rect 6683 44572 6749 44573
rect 6683 44508 6684 44572
rect 6748 44508 6749 44572
rect 6683 44507 6749 44508
rect 7235 44572 7301 44573
rect 7235 44508 7236 44572
rect 7300 44508 7301 44572
rect 7235 44507 7301 44508
rect 7787 44572 7853 44573
rect 7787 44508 7788 44572
rect 7852 44508 7853 44572
rect 7787 44507 7853 44508
rect 8339 44572 8405 44573
rect 8339 44508 8340 44572
rect 8404 44508 8405 44572
rect 8339 44507 8405 44508
rect 8891 44572 8957 44573
rect 8891 44508 8892 44572
rect 8956 44508 8957 44572
rect 8891 44507 8957 44508
rect 9443 44572 9509 44573
rect 9443 44508 9444 44572
rect 9508 44508 9509 44572
rect 9443 44507 9509 44508
rect 9995 44572 10061 44573
rect 9995 44508 9996 44572
rect 10060 44508 10061 44572
rect 9995 44507 10061 44508
rect 10547 44572 10613 44573
rect 10547 44508 10548 44572
rect 10612 44508 10613 44572
rect 10547 44507 10613 44508
rect 2912 44032 2920 44096
rect 2984 44032 3000 44096
rect 3064 44032 3080 44096
rect 3144 44032 3160 44096
rect 3224 44032 3232 44096
rect 2912 43008 3232 44032
rect 11102 43893 11162 45152
rect 11654 44709 11714 45152
rect 11651 44708 11717 44709
rect 11651 44644 11652 44708
rect 11716 44644 11717 44708
rect 11651 44643 11717 44644
rect 12206 44573 12266 45152
rect 12758 44573 12818 45152
rect 13310 44573 13370 45152
rect 13862 44573 13922 45152
rect 12203 44572 12269 44573
rect 12203 44508 12204 44572
rect 12268 44508 12269 44572
rect 12203 44507 12269 44508
rect 12755 44572 12821 44573
rect 12755 44508 12756 44572
rect 12820 44508 12821 44572
rect 12755 44507 12821 44508
rect 13307 44572 13373 44573
rect 13307 44508 13308 44572
rect 13372 44508 13373 44572
rect 13307 44507 13373 44508
rect 13859 44572 13925 44573
rect 13859 44508 13860 44572
rect 13924 44508 13925 44572
rect 13859 44507 13925 44508
rect 14414 43893 14474 45152
rect 14966 44709 15026 45152
rect 14963 44708 15029 44709
rect 14963 44644 14964 44708
rect 15028 44644 15029 44708
rect 14963 44643 15029 44644
rect 15518 44573 15578 45152
rect 16070 44573 16130 45152
rect 16622 44573 16682 45152
rect 17174 44573 17234 45152
rect 17726 44709 17786 45152
rect 17723 44708 17789 44709
rect 17723 44644 17724 44708
rect 17788 44644 17789 44708
rect 17723 44643 17789 44644
rect 15515 44572 15581 44573
rect 15515 44508 15516 44572
rect 15580 44508 15581 44572
rect 15515 44507 15581 44508
rect 16067 44572 16133 44573
rect 16067 44508 16068 44572
rect 16132 44508 16133 44572
rect 16067 44507 16133 44508
rect 16619 44572 16685 44573
rect 16619 44508 16620 44572
rect 16684 44508 16685 44572
rect 16619 44507 16685 44508
rect 17171 44572 17237 44573
rect 17171 44508 17172 44572
rect 17236 44508 17237 44572
rect 17171 44507 17237 44508
rect 11099 43892 11165 43893
rect 11099 43828 11100 43892
rect 11164 43828 11165 43892
rect 11099 43827 11165 43828
rect 14411 43892 14477 43893
rect 14411 43828 14412 43892
rect 14476 43828 14477 43892
rect 14411 43827 14477 43828
rect 18278 43485 18338 45152
rect 18830 43757 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 18827 43756 18893 43757
rect 18827 43692 18828 43756
rect 18892 43692 18893 43756
rect 18827 43691 18893 43692
rect 18275 43484 18341 43485
rect 18275 43420 18276 43484
rect 18340 43420 18341 43484
rect 18275 43419 18341 43420
rect 2912 42944 2920 43008
rect 2984 42944 3000 43008
rect 3064 42944 3080 43008
rect 3144 42944 3160 43008
rect 3224 42944 3232 43008
rect 2912 41920 3232 42944
rect 17907 42124 17973 42125
rect 17907 42060 17908 42124
rect 17972 42060 17973 42124
rect 17907 42059 17973 42060
rect 2912 41856 2920 41920
rect 2984 41856 3000 41920
rect 3064 41856 3080 41920
rect 3144 41856 3160 41920
rect 3224 41856 3232 41920
rect 2912 40832 3232 41856
rect 2912 40768 2920 40832
rect 2984 40768 3000 40832
rect 3064 40768 3080 40832
rect 3144 40768 3160 40832
rect 3224 40768 3232 40832
rect 2912 39744 3232 40768
rect 2912 39680 2920 39744
rect 2984 39680 3000 39744
rect 3064 39680 3080 39744
rect 3144 39680 3160 39744
rect 3224 39680 3232 39744
rect 2912 38656 3232 39680
rect 15515 39404 15581 39405
rect 15515 39340 15516 39404
rect 15580 39340 15581 39404
rect 15515 39339 15581 39340
rect 2912 38592 2920 38656
rect 2984 38592 3000 38656
rect 3064 38592 3080 38656
rect 3144 38592 3160 38656
rect 3224 38592 3232 38656
rect 2912 37568 3232 38592
rect 14411 38044 14477 38045
rect 14411 37980 14412 38044
rect 14476 37980 14477 38044
rect 14411 37979 14477 37980
rect 2912 37504 2920 37568
rect 2984 37504 3000 37568
rect 3064 37504 3080 37568
rect 3144 37504 3160 37568
rect 3224 37504 3232 37568
rect 2912 34796 3232 37504
rect 10915 37092 10981 37093
rect 10915 37028 10916 37092
rect 10980 37028 10981 37092
rect 10915 37027 10981 37028
rect 9627 36956 9693 36957
rect 9627 36892 9628 36956
rect 9692 36892 9693 36956
rect 9627 36891 9693 36892
rect 6131 36684 6197 36685
rect 6131 36620 6132 36684
rect 6196 36620 6197 36684
rect 6131 36619 6197 36620
rect 3923 36548 3989 36549
rect 3923 36484 3924 36548
rect 3988 36484 3989 36548
rect 3923 36483 3989 36484
rect 3926 35730 3986 36483
rect 4981 36004 5047 36005
rect 4981 35940 4982 36004
rect 5046 35940 5047 36004
rect 4981 35939 5047 35940
rect 3834 35670 3986 35730
rect 3834 35476 3894 35670
rect 4984 35476 5044 35939
rect 6134 35476 6194 36619
rect 7327 35732 7393 35733
rect 7327 35668 7328 35732
rect 7392 35668 7393 35732
rect 7327 35667 7393 35668
rect 8485 35732 8551 35733
rect 8485 35668 8486 35732
rect 8550 35668 8551 35732
rect 9630 35730 9690 36891
rect 10918 35730 10978 37027
rect 12019 36820 12085 36821
rect 12019 36756 12020 36820
rect 12084 36756 12085 36820
rect 12019 36755 12085 36756
rect 12022 35730 12082 36755
rect 13157 36004 13223 36005
rect 13157 35940 13158 36004
rect 13222 35940 13223 36004
rect 13157 35939 13223 35940
rect 9630 35670 9716 35730
rect 8485 35667 8551 35668
rect 7330 35476 7390 35667
rect 8488 35476 8548 35667
rect 9656 35476 9716 35670
rect 10826 35670 10978 35730
rect 11992 35670 12082 35730
rect 10826 35476 10886 35670
rect 11992 35476 12052 35670
rect 13160 35476 13220 35939
rect 14414 35910 14474 37979
rect 15518 35910 15578 39339
rect 16619 36140 16685 36141
rect 16619 36076 16620 36140
rect 16684 36076 16685 36140
rect 16619 36075 16685 36076
rect 14322 35850 14474 35910
rect 15496 35850 15578 35910
rect 16622 35910 16682 36075
rect 17910 35910 17970 42059
rect 19011 39812 19077 39813
rect 19011 39748 19012 39812
rect 19076 39748 19077 39812
rect 19011 39747 19077 39748
rect 16622 35850 16724 35910
rect 14322 35476 14382 35850
rect 15496 35476 15556 35850
rect 16664 35476 16724 35850
rect 17832 35850 17970 35910
rect 17832 35476 17892 35850
rect 19014 35476 19074 39747
rect 21403 38316 21469 38317
rect 21403 38252 21404 38316
rect 21468 38252 21469 38316
rect 21403 38251 21469 38252
rect 20115 37636 20181 37637
rect 20115 37572 20116 37636
rect 20180 37572 20181 37636
rect 20115 37571 20181 37572
rect 19563 36276 19629 36277
rect 19563 36212 19564 36276
rect 19628 36212 19629 36276
rect 19563 36211 19629 36212
rect 19566 35910 19626 36211
rect 19474 35850 19626 35910
rect 20118 35910 20178 37571
rect 21035 37092 21101 37093
rect 21035 37028 21036 37092
rect 21100 37028 21101 37092
rect 21035 37027 21101 37028
rect 21038 35910 21098 37027
rect 21406 35910 21466 38251
rect 21590 36957 21650 45152
rect 22142 41173 22202 45152
rect 22694 43213 22754 45152
rect 22691 43212 22757 43213
rect 22691 43148 22692 43212
rect 22756 43148 22757 43212
rect 22691 43147 22757 43148
rect 23246 42805 23306 45152
rect 23243 42804 23309 42805
rect 23243 42740 23244 42804
rect 23308 42740 23309 42804
rect 23243 42739 23309 42740
rect 23798 41430 23858 45152
rect 24350 44981 24410 45152
rect 24347 44980 24413 44981
rect 24347 44916 24348 44980
rect 24412 44916 24413 44980
rect 24347 44915 24413 44916
rect 24531 43212 24597 43213
rect 24531 43148 24532 43212
rect 24596 43148 24597 43212
rect 24531 43147 24597 43148
rect 23614 41370 23858 41430
rect 22139 41172 22205 41173
rect 22139 41108 22140 41172
rect 22204 41108 22205 41172
rect 22139 41107 22205 41108
rect 22507 39268 22573 39269
rect 22507 39204 22508 39268
rect 22572 39204 22573 39268
rect 22507 39203 22573 39204
rect 21587 36956 21653 36957
rect 21587 36892 21588 36956
rect 21652 36892 21653 36956
rect 21587 36891 21653 36892
rect 20118 35850 20228 35910
rect 19474 35476 19534 35850
rect 20027 35732 20093 35733
rect 20027 35668 20028 35732
rect 20092 35668 20093 35732
rect 20027 35667 20093 35668
rect 20030 35476 20090 35667
rect 20168 35476 20228 35850
rect 20970 35850 21098 35910
rect 21336 35850 21466 35910
rect 21967 35868 22033 35869
rect 20970 35476 21030 35850
rect 21195 35732 21261 35733
rect 21195 35668 21196 35732
rect 21260 35668 21261 35732
rect 21195 35667 21261 35668
rect 21198 35476 21258 35667
rect 21336 35476 21396 35850
rect 21967 35804 21968 35868
rect 22032 35804 22033 35868
rect 21967 35803 22033 35804
rect 21970 35476 22030 35803
rect 22197 35732 22263 35733
rect 22197 35668 22198 35732
rect 22262 35668 22263 35732
rect 22197 35667 22263 35668
rect 22200 35476 22260 35667
rect 22510 35476 22570 39203
rect 23614 36549 23674 41370
rect 24534 38861 24594 43147
rect 24902 41430 24962 45152
rect 25454 44845 25514 45152
rect 26006 44981 26066 45152
rect 26003 44980 26069 44981
rect 26003 44916 26004 44980
rect 26068 44916 26069 44980
rect 26003 44915 26069 44916
rect 25451 44844 25517 44845
rect 25451 44780 25452 44844
rect 25516 44780 25517 44844
rect 25451 44779 25517 44780
rect 26558 44437 26618 45152
rect 27110 44437 27170 45152
rect 27662 44709 27722 45152
rect 27659 44708 27725 44709
rect 27659 44644 27660 44708
rect 27724 44644 27725 44708
rect 27659 44643 27725 44644
rect 28214 44437 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 50992 44640 51312 44656
rect 50992 44576 51000 44640
rect 51064 44576 51080 44640
rect 51144 44576 51160 44640
rect 51224 44576 51240 44640
rect 51304 44576 51312 44640
rect 26555 44436 26621 44437
rect 26555 44372 26556 44436
rect 26620 44372 26621 44436
rect 26555 44371 26621 44372
rect 27107 44436 27173 44437
rect 27107 44372 27108 44436
rect 27172 44372 27173 44436
rect 27107 44371 27173 44372
rect 28211 44436 28277 44437
rect 28211 44372 28212 44436
rect 28276 44372 28277 44436
rect 28211 44371 28277 44372
rect 31891 43756 31957 43757
rect 31891 43692 31892 43756
rect 31956 43692 31957 43756
rect 31891 43691 31957 43692
rect 27107 43076 27173 43077
rect 27107 43012 27108 43076
rect 27172 43012 27173 43076
rect 27107 43011 27173 43012
rect 24902 41370 25146 41430
rect 24531 38860 24597 38861
rect 24531 38796 24532 38860
rect 24596 38796 24597 38860
rect 24531 38795 24597 38796
rect 24899 38044 24965 38045
rect 24899 37980 24900 38044
rect 24964 37980 24965 38044
rect 24899 37979 24965 37980
rect 23795 36956 23861 36957
rect 23795 36892 23796 36956
rect 23860 36892 23861 36956
rect 23795 36891 23861 36892
rect 23611 36548 23677 36549
rect 23611 36484 23612 36548
rect 23676 36484 23677 36548
rect 23611 36483 23677 36484
rect 23531 35868 23597 35869
rect 23531 35804 23532 35868
rect 23596 35804 23597 35868
rect 23798 35866 23858 36891
rect 23531 35803 23597 35804
rect 23672 35806 23858 35866
rect 24473 35868 24539 35869
rect 22967 35732 23033 35733
rect 22967 35668 22968 35732
rect 23032 35668 23033 35732
rect 22967 35667 23033 35668
rect 23197 35732 23263 35733
rect 23197 35668 23198 35732
rect 23262 35668 23263 35732
rect 23197 35667 23263 35668
rect 22970 35476 23030 35667
rect 23200 35476 23260 35667
rect 23534 35476 23594 35803
rect 23672 35476 23732 35806
rect 24473 35804 24474 35868
rect 24538 35804 24539 35868
rect 24715 35868 24781 35869
rect 24715 35866 24716 35868
rect 24473 35803 24539 35804
rect 24694 35804 24716 35866
rect 24780 35804 24781 35868
rect 24694 35803 24781 35804
rect 24476 35476 24536 35803
rect 24694 35476 24754 35803
rect 24902 35730 24962 37979
rect 25086 36413 25146 41370
rect 26739 41308 26805 41309
rect 26739 41244 26740 41308
rect 26804 41244 26805 41308
rect 26739 41243 26805 41244
rect 26003 39540 26069 39541
rect 26003 39476 26004 39540
rect 26068 39476 26069 39540
rect 26003 39475 26069 39476
rect 25083 36412 25149 36413
rect 25083 36348 25084 36412
rect 25148 36348 25149 36412
rect 25083 36347 25149 36348
rect 25867 35868 25933 35869
rect 25867 35804 25868 35868
rect 25932 35804 25933 35868
rect 25867 35803 25933 35804
rect 24840 35670 24962 35730
rect 25209 35732 25275 35733
rect 24840 35476 24900 35670
rect 25209 35668 25210 35732
rect 25274 35668 25275 35732
rect 25209 35667 25275 35668
rect 25212 35476 25272 35667
rect 25870 35476 25930 35803
rect 26006 35476 26066 39475
rect 26473 36004 26539 36005
rect 26473 35940 26474 36004
rect 26538 35940 26539 36004
rect 26473 35939 26539 35940
rect 26476 35476 26536 35939
rect 26742 35866 26802 41243
rect 27110 35866 27170 43011
rect 28947 42804 29013 42805
rect 28947 42740 28948 42804
rect 29012 42740 29013 42804
rect 28947 42739 29013 42740
rect 27843 42396 27909 42397
rect 27843 42332 27844 42396
rect 27908 42332 27909 42396
rect 27843 42331 27909 42332
rect 27291 39132 27357 39133
rect 27291 39068 27292 39132
rect 27356 39068 27357 39132
rect 27291 39067 27357 39068
rect 26694 35806 26802 35866
rect 27038 35806 27170 35866
rect 26694 35476 26754 35806
rect 27038 35476 27098 35806
rect 27294 35730 27354 39067
rect 27475 38860 27541 38861
rect 27475 38796 27476 38860
rect 27540 38796 27541 38860
rect 27475 38795 27541 38796
rect 27478 37909 27538 38795
rect 27475 37908 27541 37909
rect 27475 37844 27476 37908
rect 27540 37844 27541 37908
rect 27475 37843 27541 37844
rect 27846 35866 27906 42331
rect 28211 42260 28277 42261
rect 28211 42196 28212 42260
rect 28276 42196 28277 42260
rect 28211 42195 28277 42196
rect 27176 35670 27354 35730
rect 27694 35806 27906 35866
rect 27176 35476 27236 35670
rect 27694 35476 27754 35806
rect 28214 35476 28274 42195
rect 28950 41037 29010 42739
rect 30971 41988 31037 41989
rect 30971 41924 30972 41988
rect 31036 41924 31037 41988
rect 30971 41923 31037 41924
rect 28947 41036 29013 41037
rect 28947 40972 28948 41036
rect 29012 40972 29013 41036
rect 28947 40971 29013 40972
rect 28947 39404 29013 39405
rect 28947 39340 28948 39404
rect 29012 39340 29013 39404
rect 28947 39339 29013 39340
rect 28395 38724 28461 38725
rect 28395 38660 28396 38724
rect 28460 38660 28461 38724
rect 28395 38659 28461 38660
rect 28398 35866 28458 38659
rect 28344 35806 28458 35866
rect 28344 35476 28404 35806
rect 28950 35476 29010 39339
rect 30235 37908 30301 37909
rect 30235 37844 30236 37908
rect 30300 37906 30301 37908
rect 30300 37846 30666 37906
rect 30300 37844 30301 37846
rect 30235 37843 30301 37844
rect 29315 37500 29381 37501
rect 29315 37436 29316 37500
rect 29380 37436 29381 37500
rect 29315 37435 29381 37436
rect 29318 35730 29378 37435
rect 30606 36821 30666 37846
rect 30603 36820 30669 36821
rect 30603 36756 30604 36820
rect 30668 36756 30669 36820
rect 30603 36755 30669 36756
rect 29509 35868 29575 35869
rect 29509 35804 29510 35868
rect 29574 35804 29575 35868
rect 29509 35803 29575 35804
rect 30197 35868 30263 35869
rect 30197 35804 30198 35868
rect 30262 35804 30263 35868
rect 30197 35803 30263 35804
rect 30695 35868 30761 35869
rect 30695 35804 30696 35868
rect 30760 35804 30761 35868
rect 30974 35866 31034 41923
rect 31894 39813 31954 43691
rect 50992 43552 51312 44576
rect 50992 43488 51000 43552
rect 51064 43488 51080 43552
rect 51144 43488 51160 43552
rect 51224 43488 51240 43552
rect 51304 43488 51312 43552
rect 50992 42464 51312 43488
rect 50992 42400 51000 42464
rect 51064 42400 51080 42464
rect 51144 42400 51160 42464
rect 51224 42400 51240 42464
rect 51304 42400 51312 42464
rect 36123 41716 36189 41717
rect 36123 41652 36124 41716
rect 36188 41652 36189 41716
rect 36123 41651 36189 41652
rect 35019 41444 35085 41445
rect 35019 41380 35020 41444
rect 35084 41380 35085 41444
rect 35019 41379 35085 41380
rect 32995 40900 33061 40901
rect 32995 40836 32996 40900
rect 33060 40836 33061 40900
rect 32995 40835 33061 40836
rect 32075 40084 32141 40085
rect 32075 40020 32076 40084
rect 32140 40020 32141 40084
rect 32075 40019 32141 40020
rect 31891 39812 31957 39813
rect 31891 39748 31892 39812
rect 31956 39748 31957 39812
rect 31891 39747 31957 39748
rect 31339 39540 31405 39541
rect 31339 39476 31340 39540
rect 31404 39476 31405 39540
rect 31339 39475 31405 39476
rect 31342 35866 31402 39475
rect 32078 38450 32138 40019
rect 31894 38390 32138 38450
rect 31894 36410 31954 38390
rect 32998 38317 33058 40835
rect 32995 38316 33061 38317
rect 32995 38252 32996 38316
rect 33060 38252 33061 38316
rect 32995 38251 33061 38252
rect 32075 37908 32141 37909
rect 32075 37844 32076 37908
rect 32140 37844 32141 37908
rect 32075 37843 32141 37844
rect 32995 37908 33061 37909
rect 32995 37844 32996 37908
rect 33060 37844 33061 37908
rect 32995 37843 33061 37844
rect 32078 37365 32138 37843
rect 32075 37364 32141 37365
rect 32075 37300 32076 37364
rect 32140 37300 32141 37364
rect 32075 37299 32141 37300
rect 32443 37228 32509 37229
rect 32443 37164 32444 37228
rect 32508 37164 32509 37228
rect 32443 37163 32509 37164
rect 30974 35806 31101 35866
rect 30695 35803 30761 35804
rect 29200 35670 29378 35730
rect 29200 35476 29260 35670
rect 29512 35476 29572 35803
rect 29967 35732 30033 35733
rect 29967 35668 29968 35732
rect 30032 35668 30033 35732
rect 29967 35667 30033 35668
rect 29970 35476 30030 35667
rect 30200 35476 30260 35803
rect 30698 35476 30758 35803
rect 31041 35476 31101 35806
rect 31200 35806 31402 35866
rect 31710 36350 31954 36410
rect 31200 35476 31260 35806
rect 31710 35476 31770 36350
rect 31845 35868 31911 35869
rect 31845 35804 31846 35868
rect 31910 35804 31911 35868
rect 31845 35803 31911 35804
rect 31848 35476 31908 35803
rect 32446 35730 32506 37163
rect 32811 37092 32877 37093
rect 32811 37028 32812 37092
rect 32876 37028 32877 37092
rect 32811 37027 32877 37028
rect 32814 35730 32874 37027
rect 32998 35730 33058 37843
rect 33731 37364 33797 37365
rect 33731 37300 33732 37364
rect 33796 37300 33797 37364
rect 33731 37299 33797 37300
rect 33363 37228 33429 37229
rect 33363 37164 33364 37228
rect 33428 37164 33429 37228
rect 33363 37163 33429 37164
rect 33366 35730 33426 37163
rect 33734 35730 33794 37299
rect 34043 36004 34109 36005
rect 34043 35940 34044 36004
rect 34108 35940 34109 36004
rect 34043 35939 34109 35940
rect 32446 35670 32536 35730
rect 32814 35670 32938 35730
rect 32998 35670 33076 35730
rect 33366 35670 33518 35730
rect 32476 35476 32536 35670
rect 32878 35476 32938 35670
rect 33016 35476 33076 35670
rect 33458 35476 33518 35670
rect 33694 35670 33794 35730
rect 33694 35476 33754 35670
rect 34046 35476 34106 35939
rect 34181 35868 34247 35869
rect 34181 35804 34182 35868
rect 34246 35804 34247 35868
rect 34181 35803 34247 35804
rect 34184 35476 34244 35803
rect 35022 35730 35082 41379
rect 35387 38588 35453 38589
rect 35387 38524 35388 38588
rect 35452 38524 35453 38588
rect 35387 38523 35453 38524
rect 35197 35868 35263 35869
rect 35197 35804 35198 35868
rect 35262 35804 35263 35868
rect 35197 35803 35263 35804
rect 34970 35670 35082 35730
rect 34970 35476 35030 35670
rect 35200 35476 35260 35803
rect 35390 35730 35450 38523
rect 35352 35670 35450 35730
rect 36126 35730 36186 41651
rect 50992 41376 51312 42400
rect 50992 41312 51000 41376
rect 51064 41312 51080 41376
rect 51144 41312 51160 41376
rect 51224 41312 51240 41376
rect 51304 41312 51312 41376
rect 50992 40288 51312 41312
rect 50992 40224 51000 40288
rect 51064 40224 51080 40288
rect 51144 40224 51160 40288
rect 51224 40224 51240 40288
rect 51304 40224 51312 40288
rect 44587 40220 44653 40221
rect 44587 40156 44588 40220
rect 44652 40156 44653 40220
rect 44587 40155 44653 40156
rect 42379 37228 42445 37229
rect 42379 37164 42380 37228
rect 42444 37164 42445 37228
rect 42379 37163 42445 37164
rect 39987 36684 40053 36685
rect 39987 36620 39988 36684
rect 40052 36620 40053 36684
rect 39987 36619 40053 36620
rect 37685 36004 37751 36005
rect 37685 35940 37686 36004
rect 37750 35940 37751 36004
rect 37685 35939 37751 35940
rect 36517 35732 36583 35733
rect 36126 35670 36278 35730
rect 35352 35476 35412 35670
rect 36218 35476 36278 35670
rect 36517 35668 36518 35732
rect 36582 35668 36583 35732
rect 36517 35667 36583 35668
rect 36520 35476 36580 35667
rect 37688 35476 37748 35939
rect 38853 35868 38919 35869
rect 38853 35804 38854 35868
rect 38918 35804 38919 35868
rect 38853 35803 38919 35804
rect 38856 35476 38916 35803
rect 39990 35730 40050 36619
rect 41183 35732 41249 35733
rect 39990 35670 40084 35730
rect 40024 35476 40084 35670
rect 41183 35668 41184 35732
rect 41248 35668 41249 35732
rect 42382 35730 42442 37163
rect 43525 35868 43591 35869
rect 43525 35804 43526 35868
rect 43590 35804 43591 35868
rect 43525 35803 43591 35804
rect 41183 35667 41249 35668
rect 42360 35670 42442 35730
rect 41186 35476 41246 35667
rect 42360 35476 42420 35670
rect 43528 35476 43588 35803
rect 44590 35730 44650 40155
rect 46979 39812 47045 39813
rect 46979 39748 46980 39812
rect 47044 39748 47045 39812
rect 46979 39747 47045 39748
rect 45875 36820 45941 36821
rect 45875 36756 45876 36820
rect 45940 36756 45941 36820
rect 45875 36755 45941 36756
rect 44590 35670 44742 35730
rect 44682 35476 44742 35670
rect 45878 35476 45938 36755
rect 46982 35730 47042 39747
rect 50992 39200 51312 40224
rect 50992 39136 51000 39200
rect 51064 39136 51080 39200
rect 51144 39136 51160 39200
rect 51224 39136 51240 39200
rect 51304 39136 51312 39200
rect 50992 38112 51312 39136
rect 50992 38048 51000 38112
rect 51064 38048 51080 38112
rect 51144 38048 51160 38112
rect 51224 38048 51240 38112
rect 51304 38048 51312 38112
rect 50992 37024 51312 38048
rect 50992 36960 51000 37024
rect 51064 36960 51080 37024
rect 51144 36960 51160 37024
rect 51224 36960 51240 37024
rect 51304 36960 51312 37024
rect 46982 35670 47092 35730
rect 47032 35476 47092 35670
rect 50992 35492 51312 36960
rect 2912 34732 2920 34796
rect 2984 34732 3000 34796
rect 3064 34732 3080 34796
rect 3144 34732 3160 34796
rect 3224 34732 3232 34796
rect 2912 34716 3232 34732
rect 2912 34652 2920 34716
rect 2984 34652 3000 34716
rect 3064 34652 3080 34716
rect 3144 34652 3160 34716
rect 3224 34652 3232 34716
rect 2912 34636 3232 34652
rect 2912 34572 2920 34636
rect 2984 34572 3000 34636
rect 3064 34572 3080 34636
rect 3144 34572 3160 34636
rect 3224 34572 3232 34636
rect 2912 34556 3232 34572
rect 2912 34492 2920 34556
rect 2984 34492 3000 34556
rect 3064 34492 3080 34556
rect 3144 34492 3160 34556
rect 3224 34492 3232 34556
rect 2912 34210 3232 34492
rect 50992 35428 51000 35492
rect 51064 35428 51080 35492
rect 51144 35428 51160 35492
rect 51224 35428 51240 35492
rect 51304 35428 51312 35492
rect 50992 35412 51312 35428
rect 50992 35348 51000 35412
rect 51064 35348 51080 35412
rect 51144 35348 51160 35412
rect 51224 35348 51240 35412
rect 51304 35348 51312 35412
rect 50992 35332 51312 35348
rect 50992 35268 51000 35332
rect 51064 35268 51080 35332
rect 51144 35268 51160 35332
rect 51224 35268 51240 35332
rect 51304 35268 51312 35332
rect 50992 35252 51312 35268
rect 50992 35188 51000 35252
rect 51064 35188 51080 35252
rect 51144 35188 51160 35252
rect 51224 35188 51240 35252
rect 51304 35188 51312 35252
rect 50992 34142 51312 35188
rect 51912 44096 52232 44656
rect 51912 44032 51920 44096
rect 51984 44032 52000 44096
rect 52064 44032 52080 44096
rect 52144 44032 52160 44096
rect 52224 44032 52232 44096
rect 51912 43008 52232 44032
rect 51912 42944 51920 43008
rect 51984 42944 52000 43008
rect 52064 42944 52080 43008
rect 52144 42944 52160 43008
rect 52224 42944 52232 43008
rect 51912 41920 52232 42944
rect 62619 42260 62685 42261
rect 62619 42196 62620 42260
rect 62684 42196 62685 42260
rect 62619 42195 62685 42196
rect 51912 41856 51920 41920
rect 51984 41856 52000 41920
rect 52064 41856 52080 41920
rect 52144 41856 52160 41920
rect 52224 41856 52232 41920
rect 51912 40832 52232 41856
rect 51912 40768 51920 40832
rect 51984 40768 52000 40832
rect 52064 40768 52080 40832
rect 52144 40768 52160 40832
rect 52224 40768 52232 40832
rect 51912 39744 52232 40768
rect 51912 39680 51920 39744
rect 51984 39680 52000 39744
rect 52064 39680 52080 39744
rect 52144 39680 52160 39744
rect 52224 39680 52232 39744
rect 51912 38656 52232 39680
rect 51912 38592 51920 38656
rect 51984 38592 52000 38656
rect 52064 38592 52080 38656
rect 52144 38592 52160 38656
rect 52224 38592 52232 38656
rect 51912 37568 52232 38592
rect 51912 37504 51920 37568
rect 51984 37504 52000 37568
rect 52064 37504 52080 37568
rect 52144 37504 52160 37568
rect 52224 37504 52232 37568
rect 51912 34796 52232 37504
rect 56245 35732 56311 35733
rect 56245 35668 56246 35732
rect 56310 35668 56311 35732
rect 56245 35667 56311 35668
rect 56248 35476 56308 35667
rect 51912 34732 51920 34796
rect 51984 34732 52000 34796
rect 52064 34732 52080 34796
rect 52144 34732 52160 34796
rect 52224 34732 52232 34796
rect 51912 34716 52232 34732
rect 51912 34652 51920 34716
rect 51984 34652 52000 34716
rect 52064 34652 52080 34716
rect 52144 34652 52160 34716
rect 52224 34652 52232 34716
rect 51912 34636 52232 34652
rect 51912 34572 51920 34636
rect 51984 34572 52000 34636
rect 52064 34572 52080 34636
rect 52144 34572 52160 34636
rect 52224 34572 52232 34636
rect 51912 34556 52232 34572
rect 51912 34492 51920 34556
rect 51984 34492 52000 34556
rect 52064 34492 52080 34556
rect 52144 34492 52160 34556
rect 52224 34492 52232 34556
rect 51912 34142 52232 34492
rect 62622 29243 62682 42195
rect 63539 40220 63605 40221
rect 63539 40156 63540 40220
rect 63604 40156 63605 40220
rect 63539 40155 63605 40156
rect 63355 36004 63421 36005
rect 63355 35940 63356 36004
rect 63420 35940 63421 36004
rect 63355 35939 63421 35940
rect 62619 29242 62685 29243
rect 62619 29178 62620 29242
rect 62684 29178 62685 29242
rect 62619 29177 62685 29178
rect 63358 15333 63418 35939
rect 63542 34645 63602 40155
rect 64332 37024 64652 37584
rect 64332 36960 64340 37024
rect 64404 36960 64420 37024
rect 64484 36960 64500 37024
rect 64564 36960 64580 37024
rect 64644 36960 64652 37024
rect 64091 36412 64157 36413
rect 64091 36348 64092 36412
rect 64156 36348 64157 36412
rect 64091 36347 64157 36348
rect 63907 36276 63973 36277
rect 63907 36212 63908 36276
rect 63972 36212 63973 36276
rect 63907 36211 63973 36212
rect 63723 34780 63789 34781
rect 63723 34716 63724 34780
rect 63788 34716 63789 34780
rect 63723 34715 63789 34716
rect 63539 34644 63605 34645
rect 63539 34580 63540 34644
rect 63604 34580 63605 34644
rect 63539 34579 63605 34580
rect 63355 15332 63421 15333
rect 63355 15268 63356 15332
rect 63420 15268 63421 15332
rect 63355 15267 63421 15268
rect 48943 1869 49003 2038
rect 48940 1868 49006 1869
rect 48940 1804 48941 1868
rect 49005 1804 49006 1868
rect 48940 1803 49006 1804
rect 49081 1597 49141 2038
rect 49219 1869 49279 2038
rect 49216 1868 49282 1869
rect 49216 1804 49217 1868
rect 49281 1804 49282 1868
rect 49216 1803 49282 1804
rect 49374 1733 49434 2038
rect 49676 1869 49736 2038
rect 49673 1868 49739 1869
rect 49673 1804 49674 1868
rect 49738 1804 49739 1868
rect 49673 1803 49739 1804
rect 49371 1732 49437 1733
rect 49371 1668 49372 1732
rect 49436 1668 49437 1732
rect 49834 1730 49894 2038
rect 63726 2005 63786 34715
rect 63910 6085 63970 36211
rect 63907 6084 63973 6085
rect 63907 6020 63908 6084
rect 63972 6020 63973 6084
rect 63907 6019 63973 6020
rect 64094 5949 64154 36347
rect 64332 35936 64652 36960
rect 64332 35872 64340 35936
rect 64404 35872 64420 35936
rect 64484 35872 64500 35936
rect 64564 35872 64580 35936
rect 64644 35872 64652 35936
rect 64332 34848 64652 35872
rect 64332 34784 64340 34848
rect 64404 34784 64420 34848
rect 64484 34784 64500 34848
rect 64564 34784 64580 34848
rect 64644 34784 64652 34848
rect 64332 33760 64652 34784
rect 64332 33696 64340 33760
rect 64404 33696 64420 33760
rect 64484 33696 64500 33760
rect 64564 33696 64580 33760
rect 64644 33696 64652 33760
rect 64332 32672 64652 33696
rect 64332 32608 64340 32672
rect 64404 32608 64420 32672
rect 64484 32608 64500 32672
rect 64564 32608 64580 32672
rect 64644 32608 64652 32672
rect 64332 31584 64652 32608
rect 64332 31520 64340 31584
rect 64404 31520 64420 31584
rect 64484 31520 64500 31584
rect 64564 31520 64580 31584
rect 64644 31520 64652 31584
rect 64332 30496 64652 31520
rect 64332 30432 64340 30496
rect 64404 30432 64420 30496
rect 64484 30432 64500 30496
rect 64564 30432 64580 30496
rect 64644 30432 64652 30496
rect 64332 29408 64652 30432
rect 64332 29344 64340 29408
rect 64404 29344 64420 29408
rect 64484 29344 64500 29408
rect 64564 29344 64580 29408
rect 64644 29344 64652 29408
rect 64332 28320 64652 29344
rect 64332 28256 64340 28320
rect 64404 28256 64420 28320
rect 64484 28256 64500 28320
rect 64564 28256 64580 28320
rect 64644 28256 64652 28320
rect 64332 27232 64652 28256
rect 64332 27168 64340 27232
rect 64404 27168 64420 27232
rect 64484 27168 64500 27232
rect 64564 27168 64580 27232
rect 64644 27168 64652 27232
rect 64332 26144 64652 27168
rect 64332 26080 64340 26144
rect 64404 26080 64420 26144
rect 64484 26080 64500 26144
rect 64564 26080 64580 26144
rect 64644 26080 64652 26144
rect 64332 25056 64652 26080
rect 64332 24992 64340 25056
rect 64404 24992 64420 25056
rect 64484 24992 64500 25056
rect 64564 24992 64580 25056
rect 64644 24992 64652 25056
rect 64332 23968 64652 24992
rect 64332 23904 64340 23968
rect 64404 23904 64420 23968
rect 64484 23904 64500 23968
rect 64564 23904 64580 23968
rect 64644 23904 64652 23968
rect 64332 22880 64652 23904
rect 64332 22816 64340 22880
rect 64404 22816 64420 22880
rect 64484 22816 64500 22880
rect 64564 22816 64580 22880
rect 64644 22816 64652 22880
rect 64332 21792 64652 22816
rect 64332 21728 64340 21792
rect 64404 21728 64420 21792
rect 64484 21728 64500 21792
rect 64564 21728 64580 21792
rect 64644 21728 64652 21792
rect 64332 20704 64652 21728
rect 64332 20640 64340 20704
rect 64404 20640 64420 20704
rect 64484 20640 64500 20704
rect 64564 20640 64580 20704
rect 64644 20640 64652 20704
rect 64332 19616 64652 20640
rect 64332 19552 64340 19616
rect 64404 19552 64420 19616
rect 64484 19552 64500 19616
rect 64564 19552 64580 19616
rect 64644 19552 64652 19616
rect 64332 18528 64652 19552
rect 64332 18464 64340 18528
rect 64404 18464 64420 18528
rect 64484 18464 64500 18528
rect 64564 18464 64580 18528
rect 64644 18464 64652 18528
rect 64332 17440 64652 18464
rect 64332 17376 64340 17440
rect 64404 17376 64420 17440
rect 64484 17376 64500 17440
rect 64564 17376 64580 17440
rect 64644 17376 64652 17440
rect 64332 16352 64652 17376
rect 64332 16288 64340 16352
rect 64404 16288 64420 16352
rect 64484 16288 64500 16352
rect 64564 16288 64580 16352
rect 64644 16288 64652 16352
rect 64332 15264 64652 16288
rect 64332 15200 64340 15264
rect 64404 15200 64420 15264
rect 64484 15200 64500 15264
rect 64564 15200 64580 15264
rect 64644 15200 64652 15264
rect 64332 14176 64652 15200
rect 64332 14112 64340 14176
rect 64404 14112 64420 14176
rect 64484 14112 64500 14176
rect 64564 14112 64580 14176
rect 64644 14112 64652 14176
rect 64332 13088 64652 14112
rect 64332 13024 64340 13088
rect 64404 13024 64420 13088
rect 64484 13024 64500 13088
rect 64564 13024 64580 13088
rect 64644 13024 64652 13088
rect 64332 12000 64652 13024
rect 64332 11936 64340 12000
rect 64404 11936 64420 12000
rect 64484 11936 64500 12000
rect 64564 11936 64580 12000
rect 64644 11936 64652 12000
rect 64332 10912 64652 11936
rect 64332 10848 64340 10912
rect 64404 10848 64420 10912
rect 64484 10848 64500 10912
rect 64564 10848 64580 10912
rect 64644 10848 64652 10912
rect 64332 9824 64652 10848
rect 64332 9760 64340 9824
rect 64404 9760 64420 9824
rect 64484 9760 64500 9824
rect 64564 9760 64580 9824
rect 64644 9760 64652 9824
rect 64332 8736 64652 9760
rect 64332 8672 64340 8736
rect 64404 8672 64420 8736
rect 64484 8672 64500 8736
rect 64564 8672 64580 8736
rect 64644 8672 64652 8736
rect 64332 7648 64652 8672
rect 64332 7584 64340 7648
rect 64404 7584 64420 7648
rect 64484 7584 64500 7648
rect 64564 7584 64580 7648
rect 64644 7584 64652 7648
rect 64332 6560 64652 7584
rect 64332 6496 64340 6560
rect 64404 6496 64420 6560
rect 64484 6496 64500 6560
rect 64564 6496 64580 6560
rect 64644 6496 64652 6560
rect 64091 5948 64157 5949
rect 64091 5884 64092 5948
rect 64156 5884 64157 5948
rect 64091 5883 64157 5884
rect 64332 5472 64652 6496
rect 64332 5408 64340 5472
rect 64404 5408 64420 5472
rect 64484 5408 64500 5472
rect 64564 5408 64580 5472
rect 64644 5408 64652 5472
rect 64332 4384 64652 5408
rect 64332 4320 64340 4384
rect 64404 4320 64420 4384
rect 64484 4320 64500 4384
rect 64564 4320 64580 4384
rect 64644 4320 64652 4384
rect 64332 3296 64652 4320
rect 64332 3232 64340 3296
rect 64404 3232 64420 3296
rect 64484 3232 64500 3296
rect 64564 3232 64580 3296
rect 64644 3232 64652 3296
rect 64332 2208 64652 3232
rect 64332 2144 64340 2208
rect 64404 2144 64420 2208
rect 64484 2144 64500 2208
rect 64564 2144 64580 2208
rect 64644 2144 64652 2208
rect 63723 2004 63789 2005
rect 63723 1940 63724 2004
rect 63788 1940 63789 2004
rect 63723 1939 63789 1940
rect 49834 1670 49986 1730
rect 49371 1667 49437 1668
rect 49078 1596 49144 1597
rect 49078 1532 49079 1596
rect 49143 1532 49144 1596
rect 49078 1531 49144 1532
rect 49926 1325 49986 1670
rect 49923 1324 49989 1325
rect 49923 1260 49924 1324
rect 49988 1260 49989 1324
rect 49923 1259 49989 1260
rect 64332 1120 64652 2144
rect 64332 1056 64340 1120
rect 64404 1056 64420 1120
rect 64484 1056 64500 1120
rect 64564 1056 64580 1120
rect 64644 1056 64652 1120
rect 64332 496 64652 1056
rect 65252 37568 65572 37584
rect 65252 37504 65260 37568
rect 65324 37504 65340 37568
rect 65404 37504 65420 37568
rect 65484 37504 65500 37568
rect 65564 37504 65572 37568
rect 65252 36480 65572 37504
rect 65252 36416 65260 36480
rect 65324 36416 65340 36480
rect 65404 36416 65420 36480
rect 65484 36416 65500 36480
rect 65564 36416 65572 36480
rect 65252 35392 65572 36416
rect 65252 35328 65260 35392
rect 65324 35328 65340 35392
rect 65404 35328 65420 35392
rect 65484 35328 65500 35392
rect 65564 35328 65572 35392
rect 65252 34304 65572 35328
rect 65252 34240 65260 34304
rect 65324 34240 65340 34304
rect 65404 34240 65420 34304
rect 65484 34240 65500 34304
rect 65564 34240 65572 34304
rect 65252 33216 65572 34240
rect 65252 33152 65260 33216
rect 65324 33152 65340 33216
rect 65404 33152 65420 33216
rect 65484 33152 65500 33216
rect 65564 33152 65572 33216
rect 65252 32128 65572 33152
rect 65252 32064 65260 32128
rect 65324 32064 65340 32128
rect 65404 32064 65420 32128
rect 65484 32064 65500 32128
rect 65564 32064 65572 32128
rect 65252 31040 65572 32064
rect 65252 30976 65260 31040
rect 65324 30976 65340 31040
rect 65404 30976 65420 31040
rect 65484 30976 65500 31040
rect 65564 30976 65572 31040
rect 65252 29952 65572 30976
rect 65252 29888 65260 29952
rect 65324 29888 65340 29952
rect 65404 29888 65420 29952
rect 65484 29888 65500 29952
rect 65564 29888 65572 29952
rect 65252 28864 65572 29888
rect 65252 28800 65260 28864
rect 65324 28800 65340 28864
rect 65404 28800 65420 28864
rect 65484 28800 65500 28864
rect 65564 28800 65572 28864
rect 65252 27776 65572 28800
rect 65252 27712 65260 27776
rect 65324 27712 65340 27776
rect 65404 27712 65420 27776
rect 65484 27712 65500 27776
rect 65564 27712 65572 27776
rect 65252 26688 65572 27712
rect 65252 26624 65260 26688
rect 65324 26624 65340 26688
rect 65404 26624 65420 26688
rect 65484 26624 65500 26688
rect 65564 26624 65572 26688
rect 65252 25600 65572 26624
rect 65252 25536 65260 25600
rect 65324 25536 65340 25600
rect 65404 25536 65420 25600
rect 65484 25536 65500 25600
rect 65564 25536 65572 25600
rect 65252 24512 65572 25536
rect 65252 24448 65260 24512
rect 65324 24448 65340 24512
rect 65404 24448 65420 24512
rect 65484 24448 65500 24512
rect 65564 24448 65572 24512
rect 65252 23424 65572 24448
rect 65252 23360 65260 23424
rect 65324 23360 65340 23424
rect 65404 23360 65420 23424
rect 65484 23360 65500 23424
rect 65564 23360 65572 23424
rect 65252 22336 65572 23360
rect 65252 22272 65260 22336
rect 65324 22272 65340 22336
rect 65404 22272 65420 22336
rect 65484 22272 65500 22336
rect 65564 22272 65572 22336
rect 65252 21248 65572 22272
rect 65252 21184 65260 21248
rect 65324 21184 65340 21248
rect 65404 21184 65420 21248
rect 65484 21184 65500 21248
rect 65564 21184 65572 21248
rect 65252 20160 65572 21184
rect 65252 20096 65260 20160
rect 65324 20096 65340 20160
rect 65404 20096 65420 20160
rect 65484 20096 65500 20160
rect 65564 20096 65572 20160
rect 65252 19072 65572 20096
rect 65252 19008 65260 19072
rect 65324 19008 65340 19072
rect 65404 19008 65420 19072
rect 65484 19008 65500 19072
rect 65564 19008 65572 19072
rect 65252 17984 65572 19008
rect 65252 17920 65260 17984
rect 65324 17920 65340 17984
rect 65404 17920 65420 17984
rect 65484 17920 65500 17984
rect 65564 17920 65572 17984
rect 65252 16896 65572 17920
rect 65252 16832 65260 16896
rect 65324 16832 65340 16896
rect 65404 16832 65420 16896
rect 65484 16832 65500 16896
rect 65564 16832 65572 16896
rect 65252 15808 65572 16832
rect 65252 15744 65260 15808
rect 65324 15744 65340 15808
rect 65404 15744 65420 15808
rect 65484 15744 65500 15808
rect 65564 15744 65572 15808
rect 65252 14720 65572 15744
rect 65252 14656 65260 14720
rect 65324 14656 65340 14720
rect 65404 14656 65420 14720
rect 65484 14656 65500 14720
rect 65564 14656 65572 14720
rect 65252 13632 65572 14656
rect 65252 13568 65260 13632
rect 65324 13568 65340 13632
rect 65404 13568 65420 13632
rect 65484 13568 65500 13632
rect 65564 13568 65572 13632
rect 65252 12544 65572 13568
rect 65252 12480 65260 12544
rect 65324 12480 65340 12544
rect 65404 12480 65420 12544
rect 65484 12480 65500 12544
rect 65564 12480 65572 12544
rect 65252 11456 65572 12480
rect 65252 11392 65260 11456
rect 65324 11392 65340 11456
rect 65404 11392 65420 11456
rect 65484 11392 65500 11456
rect 65564 11392 65572 11456
rect 65252 10368 65572 11392
rect 65252 10304 65260 10368
rect 65324 10304 65340 10368
rect 65404 10304 65420 10368
rect 65484 10304 65500 10368
rect 65564 10304 65572 10368
rect 65252 9280 65572 10304
rect 65252 9216 65260 9280
rect 65324 9216 65340 9280
rect 65404 9216 65420 9280
rect 65484 9216 65500 9280
rect 65564 9216 65572 9280
rect 65252 8192 65572 9216
rect 65252 8128 65260 8192
rect 65324 8128 65340 8192
rect 65404 8128 65420 8192
rect 65484 8128 65500 8192
rect 65564 8128 65572 8192
rect 65252 7104 65572 8128
rect 65252 7040 65260 7104
rect 65324 7040 65340 7104
rect 65404 7040 65420 7104
rect 65484 7040 65500 7104
rect 65564 7040 65572 7104
rect 65252 6016 65572 7040
rect 65252 5952 65260 6016
rect 65324 5952 65340 6016
rect 65404 5952 65420 6016
rect 65484 5952 65500 6016
rect 65564 5952 65572 6016
rect 65252 4928 65572 5952
rect 65252 4864 65260 4928
rect 65324 4864 65340 4928
rect 65404 4864 65420 4928
rect 65484 4864 65500 4928
rect 65564 4864 65572 4928
rect 65252 3840 65572 4864
rect 65252 3776 65260 3840
rect 65324 3776 65340 3840
rect 65404 3776 65420 3840
rect 65484 3776 65500 3840
rect 65564 3776 65572 3840
rect 65252 2752 65572 3776
rect 65252 2688 65260 2752
rect 65324 2688 65340 2752
rect 65404 2688 65420 2752
rect 65484 2688 65500 2752
rect 65564 2688 65572 2752
rect 65252 1664 65572 2688
rect 65252 1600 65260 1664
rect 65324 1600 65340 1664
rect 65404 1600 65420 1664
rect 65484 1600 65500 1664
rect 65564 1600 65572 1664
rect 65252 576 65572 1600
rect 65252 512 65260 576
rect 65324 512 65340 576
rect 65404 512 65420 576
rect 65484 512 65500 576
rect 65564 512 65572 576
rect 65252 496 65572 512
use sky130_fd_sc_hd__mux2_1  _250_
timestamp 1
transform 1 0 27048 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _251_
timestamp 1
transform 1 0 26864 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _252_
timestamp 1
transform -1 0 57960 0 1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _253_
timestamp 1
transform -1 0 14352 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _254_
timestamp 1
transform 1 0 10948 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _255_
timestamp 1
transform 1 0 10212 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _256_
timestamp 1
transform 1 0 10028 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _257_
timestamp 1
transform 1 0 21252 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _258_
timestamp 1
transform 1 0 20332 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _259_
timestamp 1
transform 1 0 9476 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _260_
timestamp 1
transform 1 0 9568 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _261_
timestamp 1
transform 1 0 6900 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _262_
timestamp 1
transform -1 0 8556 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _263_
timestamp 1
transform 1 0 10396 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _264_
timestamp 1
transform 1 0 8832 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _265_
timestamp 1
transform 1 0 8740 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _266_
timestamp 1
transform 1 0 11684 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _267_
timestamp 1
transform 1 0 10304 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _268_
timestamp 1
transform 1 0 10948 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _269_
timestamp 1
transform 1 0 58880 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _270_
timestamp 1
transform 1 0 58052 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _271_
timestamp 1
transform 1 0 57224 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _272_
timestamp 1
transform -1 0 59800 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _273_
timestamp 1
transform 1 0 59892 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _274_
timestamp 1
transform 1 0 58144 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _275_
timestamp 1
transform -1 0 55844 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _276_
timestamp 1
transform 1 0 55752 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _277_
timestamp 1
transform 1 0 57316 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _278_
timestamp 1
transform 1 0 54740 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _279_
timestamp 1
transform 1 0 54004 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _280_
timestamp 1
transform -1 0 54464 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _281_
timestamp 1
transform -1 0 56396 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _282_
timestamp 1
transform 1 0 56120 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _283_
timestamp 1
transform 1 0 55292 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _284_
timestamp 1
transform 1 0 52992 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _285_
timestamp 1
transform 1 0 52716 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _286_
timestamp 1
transform 1 0 54832 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _287_
timestamp 1
transform -1 0 18768 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _288_
timestamp 1
transform 1 0 20884 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _289_
timestamp 1
transform 1 0 53544 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _290_
timestamp 1
transform 1 0 50416 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _291_
timestamp 1
transform -1 0 49496 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _292_
timestamp 1
transform 1 0 49680 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _293_
timestamp 1
transform -1 0 51060 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _294_
timestamp 1
transform 1 0 51060 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _295_
timestamp 1
transform 1 0 48668 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _296_
timestamp 1
transform -1 0 49496 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _297_
timestamp 1
transform 1 0 49036 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _298_
timestamp 1
transform 1 0 48208 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _299_
timestamp 1
transform 1 0 47012 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _300_
timestamp 1
transform 1 0 46092 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _301_
timestamp 1
transform 1 0 47012 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _302_
timestamp 1
transform -1 0 47932 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _303_
timestamp 1
transform 1 0 47840 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _304_
timestamp 1
transform 1 0 47012 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _305_
timestamp 1
transform -1 0 45908 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _306_
timestamp 1
transform 1 0 47012 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _307_
timestamp 1
transform 1 0 46276 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _308_
timestamp 1
transform -1 0 44252 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _309_
timestamp 1
transform 1 0 43516 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _310_
timestamp 1
transform 1 0 44436 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _311_
timestamp 1
transform -1 0 42688 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _312_
timestamp 1
transform 1 0 41860 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _313_
timestamp 1
transform 1 0 42504 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _314_
timestamp 1
transform 1 0 40296 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _315_
timestamp 1
transform 1 0 40204 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _316_
timestamp 1
transform 1 0 42044 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _317_
timestamp 1
transform -1 0 16008 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _318_
timestamp 1
transform 1 0 16836 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _319_
timestamp 1
transform -1 0 40112 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _320_
timestamp 1
transform 1 0 39284 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _321_
timestamp 1
transform 1 0 36800 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _322_
timestamp 1
transform 1 0 37628 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _323_
timestamp 1
transform 1 0 35604 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _324_
timestamp 1
transform 1 0 34960 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _325_
timestamp 1
transform 1 0 36708 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _326_
timestamp 1
transform 1 0 32384 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _327_
timestamp 1
transform 1 0 31280 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _328_
timestamp 1
transform 1 0 32108 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _329_
timestamp 1
transform 1 0 30820 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _330_
timestamp 1
transform 1 0 28980 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _331_
timestamp 1
transform 1 0 30360 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _332_
timestamp 1
transform 1 0 30636 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _333_
timestamp 1
transform 1 0 29440 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _334_
timestamp 1
transform 1 0 31556 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _335_
timestamp 1
transform 1 0 28888 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _336_
timestamp 1
transform 1 0 27692 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _337_
timestamp 1
transform -1 0 29624 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _338_
timestamp 1
transform 1 0 28060 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _339_
timestamp 1
transform 1 0 26404 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _340_
timestamp 1
transform 1 0 26864 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _341_
timestamp 1
transform 1 0 26404 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _342_
timestamp 1
transform 1 0 25484 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _343_
timestamp 1
transform 1 0 26404 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _344_
timestamp 1
transform 1 0 24656 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _345_
timestamp 1
transform 1 0 22908 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _346_
timestamp 1
transform 1 0 24104 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _347_
timestamp 1
transform 1 0 16376 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _348_
timestamp 1
transform 1 0 15180 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _349_
timestamp 1
transform 1 0 23828 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _350_
timestamp 1
transform 1 0 21436 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _351_
timestamp 1
transform 1 0 20240 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1
transform 1 0 21068 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1
transform 1 0 18676 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _354_
timestamp 1
transform 1 0 17112 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _355_
timestamp 1
transform 1 0 18676 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _356_
timestamp 1
transform 1 0 14812 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _357_
timestamp 1
transform 1 0 13892 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _358_
timestamp 1
transform 1 0 16100 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _359_
timestamp 1
transform 1 0 13984 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _360_
timestamp 1
transform 1 0 12604 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _361_
timestamp 1
transform -1 0 13340 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _362_
timestamp 1
transform 1 0 12880 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _363_
timestamp 1
transform 1 0 11592 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _364_
timestamp 1
transform 1 0 12052 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _365_
timestamp 1
transform 1 0 16100 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _366_
timestamp 1
transform 1 0 14444 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _367_
timestamp 1
transform 1 0 13708 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _368_
timestamp 1
transform 1 0 42780 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _369_
timestamp 1
transform 1 0 41860 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _370_
timestamp 1
transform 1 0 42044 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _371_
timestamp 1
transform -1 0 41492 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _372_
timestamp 1
transform -1 0 44804 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _373_
timestamp 1
transform 1 0 44436 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _374_
timestamp 1
transform 1 0 44436 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _375_
timestamp 1
transform 1 0 42688 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _376_
timestamp 1
transform 1 0 47012 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _377_
timestamp 1
transform 1 0 45540 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _378_
timestamp 1
transform 1 0 43516 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _379_
timestamp 1
transform 1 0 43424 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1
transform 1 0 17572 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _381_
timestamp 1
transform 1 0 17204 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _382_
timestamp 1
transform -1 0 46736 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _383_
timestamp 1
transform 1 0 46092 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _384_
timestamp 1
transform 1 0 52992 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _385_
timestamp 1
transform -1 0 52072 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _386_
timestamp 1
transform -1 0 51152 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _387_
timestamp 1
transform 1 0 50600 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _388_
timestamp 1
transform -1 0 65412 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _389_
timestamp 1
transform 1 0 64952 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _390_
timestamp 1
transform -1 0 64768 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _391_
timestamp 1
transform 1 0 63940 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _392_
timestamp 1
transform 1 0 65320 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _393_
timestamp 1
transform 1 0 64584 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _394_
timestamp 1
transform -1 0 65320 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _395_
timestamp 1
transform 1 0 64584 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _396_
timestamp 1
transform -1 0 65412 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _397_
timestamp 1
transform 1 0 65228 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _398_
timestamp 1
transform 1 0 64676 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _399_
timestamp 1
transform 1 0 64584 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _400_
timestamp 1
transform 1 0 64584 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _401_
timestamp 1
transform 1 0 64584 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _402_
timestamp 1
transform -1 0 65228 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _403_
timestamp 1
transform 1 0 64584 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _404_
timestamp 1
transform 1 0 64584 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _405_
timestamp 1
transform 1 0 64584 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _406_
timestamp 1
transform -1 0 65320 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _407_
timestamp 1
transform 1 0 65320 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _408_
timestamp 1
transform 1 0 64584 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _409_
timestamp 1
transform 1 0 64584 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _410_
timestamp 1
transform -1 0 65320 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _411_
timestamp 1
transform 1 0 64584 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _412_
timestamp 1
transform 1 0 64584 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _413_
timestamp 1
transform 1 0 64584 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _414_
timestamp 1
transform -1 0 65136 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _415_
timestamp 1
transform 1 0 64492 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _416_
timestamp 1
transform -1 0 64308 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _417_
timestamp 1
transform 1 0 63848 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _418_
timestamp 1
transform -1 0 64676 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _419_
timestamp 1
transform 1 0 64676 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _420_
timestamp 1
transform -1 0 19872 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _421_
timestamp 1
transform 1 0 19412 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _422_
timestamp 1
transform -1 0 40940 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _423_
timestamp 1
transform 1 0 40940 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _424_
timestamp 1
transform 1 0 39284 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _425_
timestamp 1
transform 1 0 37812 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _426_
timestamp 1
transform 1 0 37812 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _427_
timestamp 1
transform -1 0 37628 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _428_
timestamp 1
transform -1 0 39376 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _429_
timestamp 1
transform 1 0 38640 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _430_
timestamp 1
transform -1 0 37812 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _431_
timestamp 1
transform 1 0 37444 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _432_
timestamp 1
transform 1 0 35512 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _433_
timestamp 1
transform 1 0 34408 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _434_
timestamp 1
transform -1 0 35880 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _435_
timestamp 1
transform 1 0 35236 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _436_
timestamp 1
transform 1 0 33948 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _437_
timestamp 1
transform 1 0 32936 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _438_
timestamp 1
transform 1 0 34132 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _439_
timestamp 1
transform -1 0 33672 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _440_
timestamp 1
transform -1 0 34592 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _441_
timestamp 1
transform 1 0 34132 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _442_
timestamp 1
transform 1 0 32936 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _443_
timestamp 1
transform 1 0 32752 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _444_
timestamp 1
transform 1 0 35420 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _445_
timestamp 1
transform 1 0 34224 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _446_
timestamp 1
transform -1 0 34960 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _447_
timestamp 1
transform -1 0 35880 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _448_
timestamp 1
transform 1 0 64676 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _449_
timestamp 1
transform -1 0 64676 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _450_
timestamp 1
transform 1 0 64584 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _451_
timestamp 1
transform 1 0 64492 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _452_
timestamp 1
transform -1 0 64676 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _453_
timestamp 1
transform 1 0 64676 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _454_
timestamp 1
transform -1 0 64676 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _455_
timestamp 1
transform 1 0 64860 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _456_
timestamp 1
transform -1 0 29808 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _457_
timestamp 1
transform 1 0 28980 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _458_
timestamp 1
transform 1 0 30176 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _459_
timestamp 1
transform 1 0 29808 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _460_
timestamp 1
transform 1 0 22080 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _461_
timestamp 1
transform 1 0 21804 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _462_
timestamp 1
transform 1 0 28612 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _463_
timestamp 1
transform 1 0 27692 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _464_
timestamp 1
transform 1 0 25024 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _465_
timestamp 1
transform 1 0 24656 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _466_
timestamp 1
transform -1 0 26312 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _467_
timestamp 1
transform 1 0 26036 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _468_
timestamp 1
transform 1 0 23828 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _469_
timestamp 1
transform -1 0 23736 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _470_
timestamp 1
transform 1 0 25668 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _471_
timestamp 1
transform 1 0 24104 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _472_
timestamp 1
transform 1 0 12604 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _473_
timestamp 1
transform 1 0 12328 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _474_
timestamp 1
transform 1 0 22080 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _475_
timestamp 1
transform 1 0 21804 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _476_
timestamp 1
transform 1 0 11132 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _477_
timestamp 1
transform 1 0 8648 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _478_
timestamp 1
transform 1 0 21252 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _479_
timestamp 1
transform 1 0 19412 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _480_
timestamp 1
transform 1 0 51244 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _481_
timestamp 1
transform 1 0 50232 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _482_
timestamp 1
transform 1 0 17848 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _483_
timestamp 1
transform 1 0 16836 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _484_
timestamp 1
transform 1 0 39284 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _485_
timestamp 1
transform 1 0 39192 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _486_
timestamp 1
transform 1 0 16284 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _487_
timestamp 1
transform 1 0 15180 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _488_
timestamp 1
transform 1 0 23828 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _489_
timestamp 1
transform 1 0 22908 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _490_
timestamp 1
transform 1 0 18676 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _491_
timestamp 1
transform 1 0 16744 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _492_
timestamp 1
transform 1 0 48208 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _493_
timestamp 1
transform -1 0 47932 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _494_
timestamp 1
transform 1 0 20240 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _495_
timestamp 1
transform 1 0 18676 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _496_
timestamp 1
transform 1 0 40204 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _497_
timestamp 1
transform 1 0 40112 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _498_
timestamp 1
transform 1 0 22264 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _499_
timestamp 1
transform -1 0 22080 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _500_
timestamp 1
transform 1 0 26404 0 -1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _501_
timestamp 1
transform -1 0 14444 0 -1 40800
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _502_
timestamp 1
transform 1 0 8372 0 1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _503_
timestamp 1
transform 1 0 9384 0 1 40800
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _504_
timestamp 1
transform 1 0 19964 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _505_
timestamp 1
transform 1 0 8740 0 -1 40800
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _506_
timestamp 1
transform 1 0 6440 0 1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _507_
timestamp 1
transform 1 0 8556 0 -1 38624
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _508_
timestamp 1
transform 1 0 6440 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _509_
timestamp 1
transform 1 0 8464 0 -1 37536
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _510_
timestamp 1
transform -1 0 10488 0 -1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _511_
timestamp 1
transform 1 0 10028 0 1 38624
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _512_
timestamp 1
transform 1 0 57040 0 1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _513_
timestamp 1
transform 1 0 57316 0 -1 39712
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _514_
timestamp 1
transform -1 0 59800 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _515_
timestamp 1
transform 1 0 57776 0 -1 38624
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _516_
timestamp 1
transform 1 0 55200 0 -1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _517_
timestamp 1
transform -1 0 57960 0 1 37536
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _518_
timestamp 1
transform 1 0 52440 0 1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _519_
timestamp 1
transform -1 0 55200 0 -1 38624
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _520_
timestamp 1
transform -1 0 56488 0 -1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _521_
timestamp 1
transform 1 0 54924 0 -1 40800
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _522_
timestamp 1
transform 1 0 52164 0 -1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _523_
timestamp 1
transform -1 0 54924 0 -1 40800
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _524_
timestamp 1
transform -1 0 20884 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _525_
timestamp 1
transform -1 0 52716 0 1 41888
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _526_
timestamp 1
transform -1 0 51428 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _527_
timestamp 1
transform 1 0 49128 0 -1 40800
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _528_
timestamp 1
transform -1 0 50232 0 -1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _529_
timestamp 1
transform 1 0 48668 0 -1 38624
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _530_
timestamp 1
transform -1 0 49496 0 1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _531_
timestamp 1
transform 1 0 47380 0 1 41888
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _532_
timestamp 1
transform 1 0 45080 0 -1 44064
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _533_
timestamp 1
transform -1 0 47656 0 1 42976
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _534_
timestamp 1
transform 1 0 45080 0 -1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _535_
timestamp 1
transform -1 0 47380 0 1 41888
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _536_
timestamp 1
transform 1 0 44896 0 -1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _537_
timestamp 1
transform -1 0 47012 0 1 39712
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _538_
timestamp 1
transform 1 0 43056 0 -1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _539_
timestamp 1
transform -1 0 45356 0 -1 38624
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _540_
timestamp 1
transform 1 0 40848 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _541_
timestamp 1
transform -1 0 43332 0 1 38624
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _542_
timestamp 1
transform 1 0 39560 0 -1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _543_
timestamp 1
transform -1 0 42044 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _544_
timestamp 1
transform 1 0 14168 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _545_
timestamp 1
transform -1 0 40204 0 -1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _546_
timestamp 1
transform 1 0 36708 0 -1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _547_
timestamp 1
transform 1 0 37168 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _548_
timestamp 1
transform 1 0 34776 0 -1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _549_
timestamp 1
transform -1 0 37168 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _550_
timestamp 1
transform 1 0 29624 0 -1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _551_
timestamp 1
transform 1 0 31924 0 -1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _552_
timestamp 1
transform 1 0 28520 0 -1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _553_
timestamp 1
transform 1 0 29808 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _554_
timestamp 1
transform 1 0 29348 0 -1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _555_
timestamp 1
transform -1 0 32108 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _556_
timestamp 1
transform 1 0 27048 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _557_
timestamp 1
transform 1 0 28980 0 1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _558_
timestamp 1
transform 1 0 24380 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _559_
timestamp 1
transform 1 0 26220 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _560_
timestamp 1
transform 1 0 24472 0 -1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _561_
timestamp 1
transform -1 0 27048 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _562_
timestamp 1
transform 1 0 22448 0 -1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _563_
timestamp 1
transform 1 0 23644 0 -1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _564_
timestamp 1
transform 1 0 14720 0 1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _565_
timestamp 1
transform 1 0 23368 0 -1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _566_
timestamp 1
transform 1 0 19320 0 -1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _567_
timestamp 1
transform 1 0 20516 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _568_
timestamp 1
transform 1 0 16560 0 -1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _569_
timestamp 1
transform 1 0 17388 0 -1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _570_
timestamp 1
transform 1 0 13524 0 -1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _571_
timestamp 1
transform -1 0 16100 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _572_
timestamp 1
transform 1 0 12144 0 -1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _573_
timestamp 1
transform 1 0 13340 0 -1 38624
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _574_
timestamp 1
transform -1 0 11408 0 1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _575_
timestamp 1
transform 1 0 11408 0 1 42976
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _576_
timestamp 1
transform 1 0 12604 0 -1 44064
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _577_
timestamp 1
transform 1 0 13524 0 1 42976
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _578_
timestamp 1
transform 1 0 40940 0 1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _579_
timestamp 1
transform -1 0 41584 0 -1 44064
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _580_
timestamp 1
transform 1 0 42136 0 -1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _581_
timestamp 1
transform 1 0 42044 0 -1 44064
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _582_
timestamp 1
transform -1 0 45540 0 -1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _583_
timestamp 1
transform 1 0 42964 0 -1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _584_
timestamp 1
transform 1 0 16192 0 1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _585_
timestamp 1
transform 1 0 45908 0 1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _586_
timestamp 1
transform -1 0 53544 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _587_
timestamp 1
transform 1 0 49864 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _588_
timestamp 1
transform 1 0 63940 0 -1 33184
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _589_
timestamp 1
transform 1 0 63848 0 1 34272
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _590_
timestamp 1
transform 1 0 64032 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _591_
timestamp 1
transform 1 0 64032 0 -1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _592_
timestamp 1
transform 1 0 64032 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _593_
timestamp 1
transform 1 0 64032 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _594_
timestamp 1
transform 1 0 64032 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _595_
timestamp 1
transform 1 0 64032 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _596_
timestamp 1
transform 1 0 64032 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _597_
timestamp 1
transform 1 0 64032 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _598_
timestamp 1
transform 1 0 64032 0 -1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _599_
timestamp 1
transform 1 0 64032 0 -1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _600_
timestamp 1
transform 1 0 64032 0 -1 31008
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _601_
timestamp 1
transform 1 0 64032 0 1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _602_
timestamp 1
transform 1 0 63112 0 -1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _603_
timestamp 1
transform 1 0 63848 0 -1 36448
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _604_
timestamp 1
transform 1 0 18400 0 -1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _605_
timestamp 1
transform 1 0 40388 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _606_
timestamp 1
transform 1 0 37168 0 1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _607_
timestamp 1
transform 1 0 37352 0 -1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _608_
timestamp 1
transform -1 0 38548 0 -1 44064
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _609_
timestamp 1
transform 1 0 37168 0 1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _610_
timestamp 1
transform 1 0 33672 0 -1 44064
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _611_
timestamp 1
transform 1 0 34868 0 1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _612_
timestamp 1
transform 1 0 32108 0 -1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _613_
timestamp 1
transform -1 0 34040 0 1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _614_
timestamp 1
transform 1 0 32108 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _615_
timestamp 1
transform 1 0 31924 0 -1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _616_
timestamp 1
transform 1 0 33212 0 -1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _617_
timestamp 1
transform -1 0 35972 0 1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _618_
timestamp 1
transform 1 0 64032 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _619_
timestamp 1
transform 1 0 64032 0 -1 12512
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _620_
timestamp 1
transform 1 0 63848 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _621_
timestamp 1
transform 1 0 63848 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _622_
timestamp 1
transform 1 0 27508 0 -1 44064
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _623_
timestamp 1
transform 1 0 29348 0 -1 44064
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _624_
timestamp 1
transform 1 0 21252 0 -1 44064
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _625_
timestamp 1
transform 1 0 26864 0 1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _626_
timestamp 1
transform 1 0 24196 0 1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _627_
timestamp 1
transform -1 0 26312 0 -1 44064
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _628_
timestamp 1
transform 1 0 23828 0 -1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _629_
timestamp 1
transform 1 0 23092 0 -1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _630_
timestamp 1
transform 1 0 11592 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _631_
timestamp 1
transform 1 0 21252 0 -1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _632_
timestamp 1
transform 1 0 7912 0 -1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _633_
timestamp 1
transform 1 0 19044 0 -1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _634_
timestamp 1
transform 1 0 49956 0 -1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _635_
timestamp 1
transform 1 0 16008 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _636_
timestamp 1
transform 1 0 37352 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _637_
timestamp 1
transform 1 0 14996 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _638_
timestamp 1
transform 1 0 21528 0 -1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _639_
timestamp 1
transform 1 0 16100 0 -1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _640_
timestamp 1
transform -1 0 48208 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _641_
timestamp 1
transform -1 0 19412 0 -1 44064
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _642_
timestamp 1
transform 1 0 39284 0 -1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _643_
timestamp 1
transform -1 0 21712 0 1 42976
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  _666_
timestamp 1
transform 1 0 15640 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _667_
timestamp 1
transform -1 0 19044 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1
transform -1 0 22264 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1
transform 1 0 22264 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1
transform -1 0 30360 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1
transform -1 0 64032 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1
transform -1 0 64768 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1
transform -1 0 35144 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1
transform 1 0 32936 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1
transform 1 0 34868 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1
transform 1 0 35052 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1
transform 1 0 36800 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1
transform 1 0 36984 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1
transform -1 0 37812 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1
transform -1 0 64676 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1
transform -1 0 64676 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1
transform -1 0 64584 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1
transform 1 0 64400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1
transform -1 0 64860 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1
transform -1 0 64676 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1
transform -1 0 64952 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1
transform -1 0 64124 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1
transform 1 0 50140 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1
transform -1 0 19688 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1
transform -1 0 43516 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1
transform -1 0 45448 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1
transform -1 0 42044 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1
transform -1 0 16284 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1
transform -1 0 17848 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1
transform 1 0 17848 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1
transform -1 0 25668 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1
transform -1 0 35420 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1
transform -1 0 52992 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1
transform 1 0 50232 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1
transform 1 0 55568 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1
transform 1 0 55384 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ui_in[3]
timestamp 1
transform 1 0 35328 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ui_in[4]
timestamp 1
transform 1 0 36708 0 -1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_ui_in[3]
timestamp 1
transform -1 0 27048 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_ui_in[4]
timestamp 1
transform 1 0 27048 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_ui_in[3]
timestamp 1
transform -1 0 37628 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_ui_in[4]
timestamp 1
transform -1 0 39468 0 -1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_ui_in[3]
timestamp 1
transform -1 0 18584 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_ui_in[4]
timestamp 1
transform -1 0 18584 0 1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_ui_in[3]
timestamp 1
transform 1 0 18768 0 -1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_ui_in[4]
timestamp 1
transform -1 0 21896 0 1 41888
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_ui_in[3]
timestamp 1
transform 1 0 54924 0 -1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_ui_in[4]
timestamp 1
transform 1 0 64124 0 -1 32096
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_ui_in[3]
timestamp 1
transform 1 0 63848 0 1 23392
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_ui_in[4]
timestamp 1
transform 1 0 63848 0 1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_ui_in[3]
timestamp 1
transform -1 0 46276 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_ui_in[4]
timestamp 1
transform 1 0 41860 0 -1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_ui_in[3]
timestamp 1
transform 1 0 52164 0 -1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_ui_in[4]
timestamp 1
transform 1 0 51152 0 1 40800
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinvlp_4  clkload0
timestamp 1
transform 1 0 25668 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__clkinvlp_4  clkload1
timestamp 1
transform 1 0 36064 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  clkload2
timestamp 1
transform 1 0 17020 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__inv_6  clkload3
timestamp 1
transform 1 0 54004 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  clkload4
timestamp 1
transform 1 0 63848 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_8  clkload5
timestamp 1
transform 1 0 43332 0 1 40800
box -38 -48 1050 592
use sky130_fd_sc_hd__bufinv_16  clkload6
timestamp 1
transform 1 0 51796 0 1 39712
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_2  clkload7
timestamp 1
transform 1 0 27232 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__clkinvlp_4  clkload8
timestamp 1
transform 1 0 38640 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  clkload9
timestamp 1
transform 1 0 16100 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__clkinvlp_4  clkload10
timestamp 1
transform -1 0 57040 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__clkinvlp_4  clkload11
timestamp 1
transform -1 0 64400 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  clkload12
timestamp 1
transform 1 0 41400 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  clkload13
timestamp 1
transform 1 0 51060 0 -1 41888
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout5
timestamp 1
transform -1 0 14444 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout6
timestamp 1
transform 1 0 31556 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout7
timestamp 1
transform 1 0 54740 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout8
timestamp 1
transform 1 0 56948 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout9
timestamp 1
transform -1 0 17480 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout10
timestamp 1
transform -1 0 23644 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout11
timestamp 1
transform -1 0 24196 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout12
timestamp 1
transform -1 0 26220 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout13
timestamp 1
transform 1 0 30084 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout14
timestamp 1
transform 1 0 34960 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout15
timestamp 1
transform 1 0 33672 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout16
timestamp 1
transform -1 0 29348 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout17
timestamp 1
transform 1 0 63848 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout18
timestamp 1
transform -1 0 40572 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout19
timestamp 1
transform -1 0 48392 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout20
timestamp 1
transform -1 0 40572 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout21
timestamp 1
transform -1 0 57868 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout22
timestamp 1
transform 1 0 52440 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout23
timestamp 1
transform 1 0 40388 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout24
timestamp 1
transform -1 0 21804 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout25
timestamp 1
transform -1 0 24196 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout26
timestamp 1
transform -1 0 14628 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout27
timestamp 1
transform -1 0 31740 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout28
timestamp 1
transform 1 0 30084 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp 1
transform -1 0 28888 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout30
timestamp 1
transform -1 0 65228 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout31
timestamp 1
transform 1 0 39836 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout32
timestamp 1
transform 1 0 39376 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout33
timestamp 1
transform 1 0 47748 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout34
timestamp 1
transform -1 0 54372 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout35
timestamp 1
transform -1 0 55108 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout36
timestamp 1
transform 1 0 36892 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout37
timestamp 1
transform -1 0 12236 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout38
timestamp 1
transform -1 0 14904 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout39
timestamp 1
transform -1 0 15272 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout40
timestamp 1
transform -1 0 17848 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout41
timestamp 1
transform 1 0 21712 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 1
transform -1 0 30912 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout43
timestamp 1
transform -1 0 31372 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout44
timestamp 1
transform 1 0 30636 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout45
timestamp 1
transform -1 0 31924 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout46
timestamp 1
transform 1 0 65412 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout47
timestamp 1
transform -1 0 39836 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout48
timestamp 1
transform -1 0 40940 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout49
timestamp 1
transform 1 0 46368 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout50
timestamp 1
transform 1 0 42872 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout51
timestamp 1
transform 1 0 54004 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout52
timestamp 1
transform -1 0 52532 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout53
timestamp 1
transform 1 0 52164 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout54
timestamp 1
transform 1 0 40940 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout55
timestamp 1
transform 1 0 30636 0 1 44064
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_688
timestamp 1636968456
transform 1 0 63848 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_700
timestamp 1
transform 1 0 64952 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_704
timestamp 1
transform 1 0 65320 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_688
timestamp 1
transform 1 0 63848 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_698
timestamp 1
transform 1 0 64768 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_704
timestamp 1
transform 1 0 65320 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_688
timestamp 1
transform 1 0 63848 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_706
timestamp 1
transform 1 0 65504 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_712
timestamp 1
transform 1 0 66056 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_710
timestamp 1
transform 1 0 65872 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_706
timestamp 1
transform 1 0 65504 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_712
timestamp 1
transform 1 0 66056 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_708
timestamp 1
transform 1 0 65688 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_712
timestamp 1
transform 1 0 66056 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_688
timestamp 1
transform 1 0 63848 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_710
timestamp 1
transform 1 0 65872 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_708
timestamp 1
transform 1 0 65688 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_712
timestamp 1
transform 1 0 66056 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_708
timestamp 1
transform 1 0 65688 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_712
timestamp 1
transform 1 0 66056 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_688
timestamp 1
transform 1 0 63848 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_696
timestamp 1
transform 1 0 64584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_706
timestamp 1
transform 1 0 65504 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_712
timestamp 1
transform 1 0 66056 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_712
timestamp 1
transform 1 0 66056 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_688
timestamp 1
transform 1 0 63848 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_688
timestamp 1
transform 1 0 63848 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_710
timestamp 1
transform 1 0 65872 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_688
timestamp 1
transform 1 0 63848 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_688
timestamp 1
transform 1 0 63848 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_710
timestamp 1
transform 1 0 65872 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_688
timestamp 1636968456
transform 1 0 63848 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_700
timestamp 1
transform 1 0 64952 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_704
timestamp 1
transform 1 0 65320 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_688
timestamp 1
transform 1 0 63848 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_705
timestamp 1
transform 1 0 65412 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_688
timestamp 1
transform 1 0 63848 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_705
timestamp 1
transform 1 0 65412 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_688
timestamp 1
transform 1 0 63848 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_694
timestamp 1
transform 1 0 64400 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_704
timestamp 1
transform 1 0 65320 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_712
timestamp 1
transform 1 0 66056 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_688
timestamp 1
transform 1 0 63848 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_705
timestamp 1
transform 1 0 65412 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_688
timestamp 1
transform 1 0 63848 0 -1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_688
timestamp 1636968456
transform 1 0 63848 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_700
timestamp 1
transform 1 0 64952 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_704
timestamp 1
transform 1 0 65320 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_688
timestamp 1
transform 1 0 63848 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_710
timestamp 1
transform 1 0 65872 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_688
timestamp 1636968456
transform 1 0 63848 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_700
timestamp 1636968456
transform 1 0 64952 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_712
timestamp 1
transform 1 0 66056 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_688
timestamp 1636968456
transform 1 0 63848 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_700
timestamp 1636968456
transform 1 0 64952 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_712
timestamp 1
transform 1 0 66056 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_688
timestamp 1
transform 1 0 63848 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_710
timestamp 1
transform 1 0 65872 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_688
timestamp 1
transform 1 0 63848 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_694
timestamp 1
transform 1 0 64400 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_697
timestamp 1636968456
transform 1 0 64676 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_709
timestamp 1
transform 1 0 65780 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_688
timestamp 1
transform 1 0 63848 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_694
timestamp 1
transform 1 0 64400 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_688
timestamp 1636968456
transform 1 0 63848 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_700
timestamp 1
transform 1 0 64952 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_704
timestamp 1
transform 1 0 65320 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_688
timestamp 1
transform 1 0 63848 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_694
timestamp 1
transform 1 0 64400 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_697
timestamp 1636968456
transform 1 0 64676 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_709
timestamp 1
transform 1 0 65780 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_688
timestamp 1
transform 1 0 63848 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_694
timestamp 1
transform 1 0 64400 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_688
timestamp 1
transform 1 0 63848 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_710
timestamp 1
transform 1 0 65872 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_688
timestamp 1
transform 1 0 63848 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_688
timestamp 1
transform 1 0 63848 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_688
timestamp 1
transform 1 0 63848 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_710
timestamp 1
transform 1 0 65872 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_688
timestamp 1
transform 1 0 63848 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_705
timestamp 1
transform 1 0 65412 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_688
timestamp 1
transform 1 0 63848 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_711
timestamp 1
transform 1 0 65964 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_688
timestamp 1
transform 1 0 63848 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_696
timestamp 1
transform 1 0 64584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_703
timestamp 1
transform 1 0 65228 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_688
timestamp 1
transform 1 0 63848 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_710
timestamp 1
transform 1 0 65872 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_688
timestamp 1
transform 1 0 63848 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_694
timestamp 1
transform 1 0 64400 0 1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_697
timestamp 1636968456
transform 1 0 64676 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_709
timestamp 1
transform 1 0 65780 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_704
timestamp 1
transform 1 0 65320 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_712
timestamp 1
transform 1 0 66056 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_708
timestamp 1
transform 1 0 65688 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_712
timestamp 1
transform 1 0 66056 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_688
timestamp 1
transform 1 0 63848 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_710
timestamp 1
transform 1 0 65872 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_708
timestamp 1
transform 1 0 65688 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_712
timestamp 1
transform 1 0 66056 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_694
timestamp 1
transform 1 0 64400 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_688
timestamp 1
transform 1 0 63848 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_688
timestamp 1
transform 1 0 63848 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_710
timestamp 1
transform 1 0 65872 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_688
timestamp 1
transform 1 0 63848 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_705
timestamp 1
transform 1 0 65412 0 1 26656
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_688
timestamp 1636968456
transform 1 0 63848 0 -1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_700
timestamp 1636968456
transform 1 0 64952 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_712
timestamp 1
transform 1 0 66056 0 -1 27744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_688
timestamp 1636968456
transform 1 0 63848 0 1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_700
timestamp 1636968456
transform 1 0 64952 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_712
timestamp 1
transform 1 0 66056 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_688
timestamp 1
transform 1 0 63848 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_692
timestamp 1
transform 1 0 64216 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_702
timestamp 1
transform 1 0 65136 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_710
timestamp 1
transform 1 0 65872 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_688
timestamp 1
transform 1 0 63848 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_710
timestamp 1
transform 1 0 65872 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_688
timestamp 1
transform 1 0 63848 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_694
timestamp 1
transform 1 0 64400 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_704
timestamp 1
transform 1 0 65320 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_688
timestamp 1
transform 1 0 63848 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_688
timestamp 1
transform 1 0 63848 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_710
timestamp 1
transform 1 0 65872 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_688
timestamp 1
transform 1 0 63848 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_56_705
timestamp 1
transform 1 0 65412 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_688
timestamp 1
transform 1 0 63848 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_711
timestamp 1
transform 1 0 65964 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_688
timestamp 1
transform 1 0 63848 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_709
timestamp 1
transform 1 0 65780 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_688
timestamp 1
transform 1 0 63848 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_709
timestamp 1
transform 1 0 65780 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_688
timestamp 1
transform 1 0 63848 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_688
timestamp 1
transform 1 0 63848 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_698
timestamp 1
transform 1 0 64768 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_709
timestamp 1
transform 1 0 65780 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_708
timestamp 1
transform 1 0 65688 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_712
timestamp 1
transform 1 0 66056 0 1 34272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_688
timestamp 1636968456
transform 1 0 63848 0 -1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_700
timestamp 1636968456
transform 1 0 64952 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_712
timestamp 1
transform 1 0 66056 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_706
timestamp 1
transform 1 0 65504 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_712
timestamp 1
transform 1 0 66056 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_708
timestamp 1
transform 1 0 65688 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_712
timestamp 1
transform 1 0 66056 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_697
timestamp 1
transform 1 0 64676 0 1 36448
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1636968456
transform 1 0 828 0 -1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1636968456
transform 1 0 1932 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_27
timestamp 1
transform 1 0 3036 0 -1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_29
timestamp 1636968456
transform 1 0 3220 0 -1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_41
timestamp 1636968456
transform 1 0 4324 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_53
timestamp 1
transform 1 0 5428 0 -1 37536
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1636968456
transform 1 0 5796 0 -1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1636968456
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_81
timestamp 1
transform 1 0 8004 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_67_85
timestamp 1
transform 1 0 8372 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_109
timestamp 1
transform 1 0 10580 0 -1 37536
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1636968456
transform 1 0 10948 0 -1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1636968456
transform 1 0 12052 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_137
timestamp 1
transform 1 0 13156 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1
transform 1 0 15364 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1
transform 1 0 15916 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_169
timestamp 1
transform 1 0 16100 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_173
timestamp 1
transform 1 0 16468 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_194
timestamp 1
transform 1 0 18400 0 -1 37536
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_206
timestamp 1636968456
transform 1 0 19504 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_218
timestamp 1
transform 1 0 20608 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_67_225
timestamp 1
transform 1 0 21252 0 -1 37536
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_236
timestamp 1636968456
transform 1 0 22264 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_248
timestamp 1
transform 1 0 23368 0 -1 37536
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_262
timestamp 1636968456
transform 1 0 24656 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_274
timestamp 1
transform 1 0 25760 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_281
timestamp 1
transform 1 0 26404 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_285
timestamp 1
transform 1 0 26772 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_303
timestamp 1
transform 1 0 28428 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_307
timestamp 1
transform 1 0 28796 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_309
timestamp 1
transform 1 0 28980 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_333
timestamp 1
transform 1 0 31188 0 -1 37536
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_346
timestamp 1636968456
transform 1 0 32384 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_358
timestamp 1
transform 1 0 33488 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_376
timestamp 1
transform 1 0 35144 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_388
timestamp 1
transform 1 0 36248 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_413
timestamp 1
transform 1 0 38548 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_419
timestamp 1
transform 1 0 39100 0 -1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1636968456
transform 1 0 41860 0 -1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1636968456
transform 1 0 42964 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_473
timestamp 1
transform 1 0 44068 0 -1 37536
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_477
timestamp 1636968456
transform 1 0 44436 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_489
timestamp 1
transform 1 0 45540 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_502
timestamp 1
transform 1 0 46736 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_505
timestamp 1
transform 1 0 47012 0 -1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_515
timestamp 1636968456
transform 1 0 47932 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_527
timestamp 1
transform 1 0 49036 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_531
timestamp 1
transform 1 0 49404 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_533
timestamp 1
transform 1 0 49588 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_550
timestamp 1
transform 1 0 51152 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_561
timestamp 1
transform 1 0 52164 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_567
timestamp 1
transform 1 0 52716 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_579
timestamp 1
transform 1 0 53820 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_589
timestamp 1
transform 1 0 54740 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_611
timestamp 1
transform 1 0 56764 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1
transform 1 0 57132 0 -1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_654
timestamp 1636968456
transform 1 0 60720 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_666
timestamp 1
transform 1 0 61824 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_67_673
timestamp 1
transform 1 0 62468 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_679
timestamp 1
transform 1 0 63020 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_709
timestamp 1
transform 1 0 65780 0 -1 37536
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1636968456
transform 1 0 828 0 1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1636968456
transform 1 0 1932 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1
transform 1 0 3036 0 1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1636968456
transform 1 0 3220 0 1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1636968456
transform 1 0 4324 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_53
timestamp 1
transform 1 0 5428 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_61
timestamp 1
transform 1 0 6164 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_85
timestamp 1
transform 1 0 8372 0 1 37536
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_116
timestamp 1636968456
transform 1 0 11224 0 1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_128
timestamp 1636968456
transform 1 0 12328 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_141
timestamp 1
transform 1 0 13524 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_175
timestamp 1
transform 1 0 16652 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_206
timestamp 1
transform 1 0 19504 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_214
timestamp 1
transform 1 0 20240 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_68_237
timestamp 1
transform 1 0 22356 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_68_253
timestamp 1
transform 1 0 23828 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_309
timestamp 1
transform 1 0 28980 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_313
timestamp 1
transform 1 0 29348 0 1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_351
timestamp 1636968456
transform 1 0 32844 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1
transform 1 0 33948 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_365
timestamp 1
transform 1 0 34132 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_375
timestamp 1
transform 1 0 35052 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_68_418
timestamp 1
transform 1 0 39008 0 1 37536
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1636968456
transform 1 0 39284 0 1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_453
timestamp 1636968456
transform 1 0 42228 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_465
timestamp 1
transform 1 0 43332 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1
transform 1 0 44252 0 1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_486
timestamp 1636968456
transform 1 0 45264 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_527
timestamp 1
transform 1 0 49036 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1
transform 1 0 49404 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_533
timestamp 1
transform 1 0 49588 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_68_576
timestamp 1
transform 1 0 53544 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_586
timestamp 1
transform 1 0 54464 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_68_589
timestamp 1
transform 1 0 54740 0 1 37536
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_653
timestamp 1636968456
transform 1 0 60628 0 1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_665
timestamp 1636968456
transform 1 0 61732 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_677
timestamp 1
transform 1 0 62836 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_683
timestamp 1
transform 1 0 63388 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_693
timestamp 1
transform 1 0 64308 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_699
timestamp 1
transform 1 0 64860 0 1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_701
timestamp 1636968456
transform 1 0 65044 0 1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1636968456
transform 1 0 828 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1636968456
transform 1 0 1932 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1636968456
transform 1 0 3036 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1636968456
transform 1 0 4140 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1
transform 1 0 5244 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1
transform 1 0 5612 0 -1 38624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1636968456
transform 1 0 5796 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_110
timestamp 1
transform 1 0 10672 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_178
timestamp 1
transform 1 0 16928 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_203
timestamp 1
transform 1 0 19228 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_225
timestamp 1
transform 1 0 21252 0 -1 38624
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_268
timestamp 1636968456
transform 1 0 25208 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_298
timestamp 1
transform 1 0 27968 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_306
timestamp 1
transform 1 0 28704 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_317
timestamp 1
transform 1 0 29716 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_345
timestamp 1
transform 1 0 32292 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_353
timestamp 1
transform 1 0 33028 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_413
timestamp 1
transform 1 0 38548 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1
transform 1 0 41124 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1
transform 1 0 41676 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_513
timestamp 1
transform 1 0 47748 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_521
timestamp 1
transform 1 0 48484 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1
transform 1 0 51428 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1
transform 1 0 51980 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_569
timestamp 1
transform 1 0 52900 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_614
timestamp 1
transform 1 0 57040 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_617
timestamp 1
transform 1 0 57316 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_621
timestamp 1
transform 1 0 57684 0 -1 38624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_645
timestamp 1636968456
transform 1 0 59892 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_657
timestamp 1636968456
transform 1 0 60996 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_669
timestamp 1
transform 1 0 62100 0 -1 38624
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_673
timestamp 1636968456
transform 1 0 62468 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_685
timestamp 1636968456
transform 1 0 63572 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_697
timestamp 1636968456
transform 1 0 64676 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_709
timestamp 1
transform 1 0 65780 0 -1 38624
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1636968456
transform 1 0 828 0 1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1636968456
transform 1 0 1932 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1
transform 1 0 3036 0 1 38624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1636968456
transform 1 0 3220 0 1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1636968456
transform 1 0 4324 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_53
timestamp 1
transform 1 0 5428 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_61
timestamp 1
transform 1 0 6164 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_85
timestamp 1
transform 1 0 8372 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_89
timestamp 1
transform 1 0 8740 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_99
timestamp 1
transform 1 0 9660 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_126
timestamp 1
transform 1 0 12144 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_130
timestamp 1
transform 1 0 12512 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_141
timestamp 1
transform 1 0 13524 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_154
timestamp 1
transform 1 0 14720 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_172
timestamp 1
transform 1 0 16376 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_240
timestamp 1
transform 1 0 22632 0 1 38624
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_287
timestamp 1636968456
transform 1 0 26956 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_299
timestamp 1
transform 1 0 28060 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1
transform 1 0 28796 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_355
timestamp 1
transform 1 0 33212 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1
transform 1 0 33948 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_385
timestamp 1
transform 1 0 35972 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_393
timestamp 1
transform 1 0 36708 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_439
timestamp 1
transform 1 0 40940 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_443
timestamp 1
transform 1 0 41308 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_465
timestamp 1
transform 1 0 43332 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_477
timestamp 1
transform 1 0 44436 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_483
timestamp 1
transform 1 0 44988 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_521
timestamp 1
transform 1 0 48484 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_533
timestamp 1
transform 1 0 49588 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_539
timestamp 1
transform 1 0 50140 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_551
timestamp 1
transform 1 0 51244 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_555
timestamp 1
transform 1 0 51612 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_584
timestamp 1
transform 1 0 54280 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_609
timestamp 1
transform 1 0 56580 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_613
timestamp 1
transform 1 0 56948 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_643
timestamp 1
transform 1 0 59708 0 1 38624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_645
timestamp 1636968456
transform 1 0 59892 0 1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_657
timestamp 1636968456
transform 1 0 60996 0 1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_669
timestamp 1636968456
transform 1 0 62100 0 1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_681
timestamp 1636968456
transform 1 0 63204 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_693
timestamp 1
transform 1 0 64308 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_699
timestamp 1
transform 1 0 64860 0 1 38624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_701
timestamp 1636968456
transform 1 0 65044 0 1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1636968456
transform 1 0 828 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1636968456
transform 1 0 1932 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1636968456
transform 1 0 3036 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1636968456
transform 1 0 4140 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1
transform 1 0 5244 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1
transform 1 0 5612 0 -1 39712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1636968456
transform 1 0 5796 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_69
timestamp 1
transform 1 0 6900 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_77
timestamp 1
transform 1 0 7636 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_87
timestamp 1
transform 1 0 8556 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_108
timestamp 1
transform 1 0 10488 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_122
timestamp 1
transform 1 0 11776 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_155
timestamp 1
transform 1 0 14812 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_218
timestamp 1
transform 1 0 20608 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_234
timestamp 1
transform 1 0 22080 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_258
timestamp 1
transform 1 0 24288 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_294
timestamp 1
transform 1 0 27600 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_333
timestamp 1
transform 1 0 31188 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_337
timestamp 1
transform 1 0 31556 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_71_369
timestamp 1
transform 1 0 34500 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_71_380
timestamp 1
transform 1 0 35512 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_390
timestamp 1
transform 1 0 36432 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_402
timestamp 1
transform 1 0 37536 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_410
timestamp 1
transform 1 0 38272 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_458
timestamp 1
transform 1 0 42688 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_502
timestamp 1
transform 1 0 46736 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_514
timestamp 1
transform 1 0 47840 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_71_558
timestamp 1
transform 1 0 51888 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_607
timestamp 1
transform 1 0 56396 0 -1 39712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_648
timestamp 1636968456
transform 1 0 60168 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_660
timestamp 1636968456
transform 1 0 61272 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_673
timestamp 1636968456
transform 1 0 62468 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_685
timestamp 1636968456
transform 1 0 63572 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_697
timestamp 1636968456
transform 1 0 64676 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_709
timestamp 1
transform 1 0 65780 0 -1 39712
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1636968456
transform 1 0 828 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1636968456
transform 1 0 1932 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1
transform 1 0 3036 0 1 39712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1636968456
transform 1 0 3220 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1636968456
transform 1 0 4324 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1636968456
transform 1 0 5428 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1636968456
transform 1 0 6532 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1
transform 1 0 7636 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1
transform 1 0 8188 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_72_85
timestamp 1
transform 1 0 8372 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_72_124
timestamp 1
transform 1 0 11960 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_130
timestamp 1
transform 1 0 12512 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_141
timestamp 1
transform 1 0 13524 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_147
timestamp 1
transform 1 0 14076 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_190
timestamp 1
transform 1 0 18032 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_197
timestamp 1
transform 1 0 18676 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_230
timestamp 1
transform 1 0 21712 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_72_253
timestamp 1
transform 1 0 23828 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_72_265
timestamp 1
transform 1 0 24932 0 1 39712
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_338
timestamp 1636968456
transform 1 0 31648 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_350
timestamp 1
transform 1 0 32752 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_354
timestamp 1
transform 1 0 33120 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_362
timestamp 1
transform 1 0 33856 0 1 39712
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1636968456
transform 1 0 34132 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_377
timestamp 1
transform 1 0 35236 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_398
timestamp 1
transform 1 0 37168 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_458
timestamp 1
transform 1 0 42688 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_464
timestamp 1
transform 1 0 43240 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_477
timestamp 1
transform 1 0 44436 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_483
timestamp 1
transform 1 0 44988 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_505
timestamp 1
transform 1 0 47012 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_514
timestamp 1
transform 1 0 47840 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_553
timestamp 1
transform 1 0 51428 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1
transform 1 0 54004 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1
transform 1 0 54556 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_589
timestamp 1
transform 1 0 54740 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_595
timestamp 1
transform 1 0 55292 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_607
timestamp 1
transform 1 0 56396 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_614
timestamp 1
transform 1 0 57040 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_634
timestamp 1
transform 1 0 58880 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_642
timestamp 1
transform 1 0 59616 0 1 39712
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_645
timestamp 1636968456
transform 1 0 59892 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_657
timestamp 1636968456
transform 1 0 60996 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_669
timestamp 1636968456
transform 1 0 62100 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_681
timestamp 1636968456
transform 1 0 63204 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_693
timestamp 1
transform 1 0 64308 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_699
timestamp 1
transform 1 0 64860 0 1 39712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_701
timestamp 1636968456
transform 1 0 65044 0 1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1636968456
transform 1 0 828 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1636968456
transform 1 0 1932 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1636968456
transform 1 0 3036 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1636968456
transform 1 0 4140 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1
transform 1 0 5244 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1
transform 1 0 5612 0 -1 40800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1636968456
transform 1 0 5796 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1636968456
transform 1 0 6900 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_81
timestamp 1
transform 1 0 8004 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_73_122
timestamp 1
transform 1 0 11776 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_73_169
timestamp 1
transform 1 0 16100 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_197
timestamp 1
transform 1 0 18676 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_73_221
timestamp 1
transform 1 0 20884 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_73_234
timestamp 1
transform 1 0 22080 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_298
timestamp 1
transform 1 0 27968 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_370
timestamp 1
transform 1 0 34592 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_393
timestamp 1
transform 1 0 36708 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_399
timestamp 1
transform 1 0 37260 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_73_429
timestamp 1
transform 1 0 40020 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_73_441
timestamp 1
transform 1 0 41124 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_73_498
timestamp 1
transform 1 0 46368 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_73_514
timestamp 1
transform 1 0 47840 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_73_561
timestamp 1
transform 1 0 52164 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_614
timestamp 1
transform 1 0 57040 0 -1 40800
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_617
timestamp 1636968456
transform 1 0 57316 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_629
timestamp 1636968456
transform 1 0 58420 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_641
timestamp 1636968456
transform 1 0 59524 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_653
timestamp 1636968456
transform 1 0 60628 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_665
timestamp 1
transform 1 0 61732 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_671
timestamp 1
transform 1 0 62284 0 -1 40800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_673
timestamp 1636968456
transform 1 0 62468 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_685
timestamp 1636968456
transform 1 0 63572 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_697
timestamp 1636968456
transform 1 0 64676 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_709
timestamp 1
transform 1 0 65780 0 -1 40800
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1636968456
transform 1 0 828 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1636968456
transform 1 0 1932 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1
transform 1 0 3036 0 1 40800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1636968456
transform 1 0 3220 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1636968456
transform 1 0 4324 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1636968456
transform 1 0 5428 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1636968456
transform 1 0 6532 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1
transform 1 0 7636 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1
transform 1 0 8188 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_85
timestamp 1
transform 1 0 8372 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_74_119
timestamp 1
transform 1 0 11500 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_150
timestamp 1
transform 1 0 14352 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_156
timestamp 1
transform 1 0 14904 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_186
timestamp 1
transform 1 0 17664 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_197
timestamp 1
transform 1 0 18676 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_240
timestamp 1
transform 1 0 22632 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_74_253
timestamp 1
transform 1 0 23828 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_74_265
timestamp 1
transform 1 0 24932 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_74_309
timestamp 1
transform 1 0 28980 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_317
timestamp 1
transform 1 0 29716 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1
transform 1 0 33948 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_430
timestamp 1
transform 1 0 40112 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_451
timestamp 1
transform 1 0 42044 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_455
timestamp 1
transform 1 0 42412 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_523
timestamp 1
transform 1 0 48668 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1
transform 1 0 49404 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_533
timestamp 1
transform 1 0 49588 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_543
timestamp 1
transform 1 0 50508 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_549
timestamp 1
transform 1 0 51060 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_585
timestamp 1
transform 1 0 54372 0 1 40800
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_624
timestamp 1636968456
transform 1 0 57960 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_636
timestamp 1
transform 1 0 59064 0 1 40800
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_74_645
timestamp 1636968456
transform 1 0 59892 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_657
timestamp 1636968456
transform 1 0 60996 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_669
timestamp 1636968456
transform 1 0 62100 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_681
timestamp 1636968456
transform 1 0 63204 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_693
timestamp 1
transform 1 0 64308 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_699
timestamp 1
transform 1 0 64860 0 1 40800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_701
timestamp 1636968456
transform 1 0 65044 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1636968456
transform 1 0 828 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1636968456
transform 1 0 1932 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1636968456
transform 1 0 3036 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1636968456
transform 1 0 4140 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1
transform 1 0 5244 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1
transform 1 0 5612 0 -1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1636968456
transform 1 0 5796 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_69
timestamp 1
transform 1 0 6900 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_77
timestamp 1
transform 1 0 7636 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_75_100
timestamp 1
transform 1 0 9752 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_75_113
timestamp 1
transform 1 0 10948 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_119
timestamp 1
transform 1 0 11500 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_151
timestamp 1
transform 1 0 14444 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_169
timestamp 1
transform 1 0 16100 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_75_198
timestamp 1
transform 1 0 18768 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1
transform 1 0 26220 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_301
timestamp 1
transform 1 0 28244 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_314
timestamp 1
transform 1 0 29440 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_320
timestamp 1
transform 1 0 29992 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_327
timestamp 1
transform 1 0 30636 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1
transform 1 0 31372 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_337
timestamp 1
transform 1 0 31556 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_361
timestamp 1
transform 1 0 33764 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_365
timestamp 1
transform 1 0 34132 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_380
timestamp 1
transform 1 0 35512 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_393
timestamp 1
transform 1 0 36708 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_423
timestamp 1
transform 1 0 39468 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_444
timestamp 1
transform 1 0 41400 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_449
timestamp 1
transform 1 0 41860 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_460
timestamp 1
transform 1 0 42872 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_75_481
timestamp 1
transform 1 0 44804 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_532
timestamp 1
transform 1 0 49496 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_587
timestamp 1
transform 1 0 54556 0 -1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_623
timestamp 1636968456
transform 1 0 57868 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_635
timestamp 1636968456
transform 1 0 58972 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_647
timestamp 1636968456
transform 1 0 60076 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_659
timestamp 1636968456
transform 1 0 61180 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_671
timestamp 1
transform 1 0 62284 0 -1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_673
timestamp 1636968456
transform 1 0 62468 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_685
timestamp 1636968456
transform 1 0 63572 0 -1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_697
timestamp 1636968456
transform 1 0 64676 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_709
timestamp 1
transform 1 0 65780 0 -1 41888
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1636968456
transform 1 0 828 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1636968456
transform 1 0 1932 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1
transform 1 0 3036 0 1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1636968456
transform 1 0 3220 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1636968456
transform 1 0 4324 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1636968456
transform 1 0 5428 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1636968456
transform 1 0 6532 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1
transform 1 0 7636 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1
transform 1 0 8188 0 1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_122
timestamp 1636968456
transform 1 0 11776 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_134
timestamp 1
transform 1 0 12880 0 1 41888
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1636968456
transform 1 0 13524 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_153
timestamp 1
transform 1 0 14628 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_174
timestamp 1
transform 1 0 16560 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_194
timestamp 1
transform 1 0 18400 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_208
timestamp 1
transform 1 0 19688 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_232
timestamp 1
transform 1 0 21896 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_238
timestamp 1
transform 1 0 22448 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_242
timestamp 1
transform 1 0 22816 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_282
timestamp 1
transform 1 0 26496 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_306
timestamp 1
transform 1 0 28704 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_317
timestamp 1
transform 1 0 29716 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_321
timestamp 1
transform 1 0 30084 0 1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_330
timestamp 1636968456
transform 1 0 30912 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_359
timestamp 1
transform 1 0 33580 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_374
timestamp 1
transform 1 0 34960 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_392
timestamp 1
transform 1 0 36616 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_418
timestamp 1
transform 1 0 39008 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_429
timestamp 1
transform 1 0 40020 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_448
timestamp 1
transform 1 0 41768 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1
transform 1 0 44252 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_533
timestamp 1
transform 1 0 49588 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_541
timestamp 1
transform 1 0 50324 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_76_585
timestamp 1
transform 1 0 54372 0 1 41888
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_593
timestamp 1636968456
transform 1 0 55108 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_605
timestamp 1636968456
transform 1 0 56212 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_617
timestamp 1636968456
transform 1 0 57316 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_629
timestamp 1636968456
transform 1 0 58420 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_641
timestamp 1
transform 1 0 59524 0 1 41888
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_645
timestamp 1636968456
transform 1 0 59892 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_657
timestamp 1636968456
transform 1 0 60996 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_669
timestamp 1636968456
transform 1 0 62100 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_681
timestamp 1636968456
transform 1 0 63204 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_693
timestamp 1
transform 1 0 64308 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_699
timestamp 1
transform 1 0 64860 0 1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_701
timestamp 1636968456
transform 1 0 65044 0 1 41888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1636968456
transform 1 0 828 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1636968456
transform 1 0 1932 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1636968456
transform 1 0 3036 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1636968456
transform 1 0 4140 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1
transform 1 0 5244 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1
transform 1 0 5612 0 -1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1636968456
transform 1 0 5796 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1636968456
transform 1 0 6900 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1636968456
transform 1 0 8004 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1636968456
transform 1 0 9108 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1
transform 1 0 10212 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1
transform 1 0 10764 0 -1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1636968456
transform 1 0 10948 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_189
timestamp 1
transform 1 0 17940 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_193
timestamp 1
transform 1 0 18308 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1
transform 1 0 21068 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_265
timestamp 1
transform 1 0 24932 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_77_284
timestamp 1
transform 1 0 26680 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_308
timestamp 1
transform 1 0 28888 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_318
timestamp 1
transform 1 0 29808 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_331
timestamp 1
transform 1 0 31004 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1
transform 1 0 31372 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_337
timestamp 1
transform 1 0 31556 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_372
timestamp 1
transform 1 0 34776 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_393
timestamp 1
transform 1 0 36708 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_435
timestamp 1
transform 1 0 40572 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_77_445
timestamp 1
transform 1 0 41492 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_77_449
timestamp 1
transform 1 0 41860 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_77_481
timestamp 1
transform 1 0 44804 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_514
timestamp 1
transform 1 0 47840 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_536
timestamp 1
transform 1 0 49864 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_77_557
timestamp 1
transform 1 0 51796 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_77_565
timestamp 1
transform 1 0 52532 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_573
timestamp 1
transform 1 0 53268 0 -1 42976
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_584
timestamp 1636968456
transform 1 0 54280 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_596
timestamp 1636968456
transform 1 0 55384 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_608
timestamp 1
transform 1 0 56488 0 -1 42976
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_77_617
timestamp 1636968456
transform 1 0 57316 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_629
timestamp 1636968456
transform 1 0 58420 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_641
timestamp 1636968456
transform 1 0 59524 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_653
timestamp 1636968456
transform 1 0 60628 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_665
timestamp 1
transform 1 0 61732 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_671
timestamp 1
transform 1 0 62284 0 -1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_673
timestamp 1636968456
transform 1 0 62468 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_685
timestamp 1636968456
transform 1 0 63572 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_697
timestamp 1636968456
transform 1 0 64676 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_709
timestamp 1
transform 1 0 65780 0 -1 42976
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1636968456
transform 1 0 828 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1636968456
transform 1 0 1932 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1
transform 1 0 3036 0 1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1636968456
transform 1 0 3220 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1636968456
transform 1 0 4324 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1636968456
transform 1 0 5428 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1636968456
transform 1 0 6532 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1
transform 1 0 7636 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1
transform 1 0 8188 0 1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1636968456
transform 1 0 8372 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_97
timestamp 1
transform 1 0 9476 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1
transform 1 0 13340 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_190
timestamp 1
transform 1 0 18032 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1
transform 1 0 23644 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_286
timestamp 1
transform 1 0 26864 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_339
timestamp 1
transform 1 0 31740 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_343
timestamp 1
transform 1 0 32108 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_393
timestamp 1
transform 1 0 36708 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_397
timestamp 1
transform 1 0 37076 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_418
timestamp 1
transform 1 0 39008 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_486
timestamp 1
transform 1 0 45264 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_490
timestamp 1
transform 1 0 45632 0 1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1636968456
transform 1 0 49588 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_545
timestamp 1
transform 1 0 50692 0 1 42976
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_565
timestamp 1636968456
transform 1 0 52532 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_577
timestamp 1
transform 1 0 53636 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_585
timestamp 1
transform 1 0 54372 0 1 42976
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1636968456
transform 1 0 54740 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1636968456
transform 1 0 55844 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_613
timestamp 1636968456
transform 1 0 56948 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_625
timestamp 1636968456
transform 1 0 58052 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_637
timestamp 1
transform 1 0 59156 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_643
timestamp 1
transform 1 0 59708 0 1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_645
timestamp 1636968456
transform 1 0 59892 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_657
timestamp 1636968456
transform 1 0 60996 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_669
timestamp 1636968456
transform 1 0 62100 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_681
timestamp 1636968456
transform 1 0 63204 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_693
timestamp 1
transform 1 0 64308 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_699
timestamp 1
transform 1 0 64860 0 1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_701
timestamp 1636968456
transform 1 0 65044 0 1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1636968456
transform 1 0 828 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1636968456
transform 1 0 1932 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1636968456
transform 1 0 3036 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1636968456
transform 1 0 4140 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1
transform 1 0 5244 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1
transform 1 0 5612 0 -1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1636968456
transform 1 0 5796 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1636968456
transform 1 0 6900 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1636968456
transform 1 0 8004 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1636968456
transform 1 0 9108 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1
transform 1 0 10212 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1
transform 1 0 10764 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_113
timestamp 1
transform 1 0 10948 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_118
timestamp 1
transform 1 0 11408 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_129
timestamp 1
transform 1 0 12420 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_163
timestamp 1
transform 1 0 15548 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_184
timestamp 1
transform 1 0 17480 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_222
timestamp 1
transform 1 0 20976 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_251
timestamp 1
transform 1 0 23644 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_341
timestamp 1
transform 1 0 31924 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_79_389
timestamp 1
transform 1 0 36340 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_446
timestamp 1
transform 1 0 41584 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_449
timestamp 1
transform 1 0 41860 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_479
timestamp 1
transform 1 0 44620 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_483
timestamp 1
transform 1 0 44988 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_520
timestamp 1
transform 1 0 48392 0 -1 44064
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_530
timestamp 1636968456
transform 1 0 49312 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_542
timestamp 1636968456
transform 1 0 50416 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_554
timestamp 1
transform 1 0 51520 0 -1 44064
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1636968456
transform 1 0 52164 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1636968456
transform 1 0 53268 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1636968456
transform 1 0 54372 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1636968456
transform 1 0 55476 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1
transform 1 0 56580 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1
transform 1 0 57132 0 -1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_617
timestamp 1636968456
transform 1 0 57316 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_629
timestamp 1636968456
transform 1 0 58420 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_641
timestamp 1636968456
transform 1 0 59524 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_653
timestamp 1636968456
transform 1 0 60628 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_665
timestamp 1
transform 1 0 61732 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_671
timestamp 1
transform 1 0 62284 0 -1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_673
timestamp 1636968456
transform 1 0 62468 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_685
timestamp 1636968456
transform 1 0 63572 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_697
timestamp 1636968456
transform 1 0 64676 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_709
timestamp 1
transform 1 0 65780 0 -1 44064
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1636968456
transform 1 0 828 0 1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1636968456
transform 1 0 1932 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1
transform 1 0 3036 0 1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1636968456
transform 1 0 3220 0 1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1636968456
transform 1 0 4324 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_53
timestamp 1
transform 1 0 5428 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_57
timestamp 1
transform 1 0 5796 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_80_64
timestamp 1
transform 1 0 6440 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_80_70
timestamp 1
transform 1 0 6992 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_80_76
timestamp 1
transform 1 0 7544 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_80_82
timestamp 1
transform 1 0 8096 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_80_88
timestamp 1
transform 1 0 8648 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_80_94
timestamp 1
transform 1 0 9200 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_80_100
timestamp 1
transform 1 0 9752 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_80_106
timestamp 1
transform 1 0 10304 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_136
timestamp 1
transform 1 0 13064 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_161
timestamp 1
transform 1 0 15364 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_169
timestamp 1
transform 1 0 16100 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_214
timestamp 1
transform 1 0 20240 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_80_240
timestamp 1
transform 1 0 22632 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1
transform 1 0 23644 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_257
timestamp 1
transform 1 0 24196 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_279
timestamp 1
transform 1 0 26220 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_335
timestamp 1
transform 1 0 31372 0 1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_337
timestamp 1636968456
transform 1 0 31556 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_349
timestamp 1
transform 1 0 32660 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_80_361
timestamp 1
transform 1 0 33764 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_80_365
timestamp 1
transform 1 0 34132 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_80_385
timestamp 1
transform 1 0 35972 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_391
timestamp 1
transform 1 0 36524 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_393
timestamp 1
transform 1 0 36708 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_418
timestamp 1
transform 1 0 39008 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_80_445
timestamp 1
transform 1 0 41492 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1
transform 1 0 44252 0 1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1636968456
transform 1 0 44436 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_489
timestamp 1
transform 1 0 45540 0 1 44064
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_519
timestamp 1636968456
transform 1 0 48300 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1
transform 1 0 49404 0 1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1636968456
transform 1 0 49588 0 1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1636968456
transform 1 0 50692 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_557
timestamp 1
transform 1 0 51796 0 1 44064
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_561
timestamp 1636968456
transform 1 0 52164 0 1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_573
timestamp 1636968456
transform 1 0 53268 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_585
timestamp 1
transform 1 0 54372 0 1 44064
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1636968456
transform 1 0 54740 0 1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1636968456
transform 1 0 55844 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_613
timestamp 1
transform 1 0 56948 0 1 44064
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_617
timestamp 1636968456
transform 1 0 57316 0 1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_629
timestamp 1636968456
transform 1 0 58420 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_641
timestamp 1
transform 1 0 59524 0 1 44064
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_645
timestamp 1636968456
transform 1 0 59892 0 1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_657
timestamp 1636968456
transform 1 0 60996 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_669
timestamp 1
transform 1 0 62100 0 1 44064
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_673
timestamp 1636968456
transform 1 0 62468 0 1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_685
timestamp 1636968456
transform 1 0 63572 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_697
timestamp 1
transform 1 0 64676 0 1 44064
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_701
timestamp 1636968456
transform 1 0 65044 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform 1 0 27416 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform 1 0 28152 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform 1 0 26680 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform -1 0 23644 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform -1 0 22908 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1
transform 1 0 24288 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1
transform -1 0 23828 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1
transform 1 0 65412 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1
transform -1 0 20332 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1
transform 1 0 32016 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1
transform 1 0 23736 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1
transform -1 0 46368 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1
transform -1 0 44252 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1
transform -1 0 66148 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1
transform -1 0 66148 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1
transform -1 0 66148 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1
transform -1 0 20240 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1
transform 1 0 15272 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1
transform 1 0 14444 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1
transform -1 0 18584 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1
transform -1 0 29716 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1
transform 1 0 32108 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1
transform 1 0 34776 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1
transform -1 0 36616 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1
transform -1 0 52440 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1
transform -1 0 66148 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1
transform -1 0 48484 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1
transform -1 0 66148 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1
transform -1 0 66148 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1
transform -1 0 66148 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1
transform 1 0 26220 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1
transform -1 0 65780 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1
transform -1 0 8556 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1
transform -1 0 30636 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1
transform -1 0 39192 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1
transform -1 0 11776 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1
transform -1 0 22632 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1
transform -1 0 47748 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1
transform -1 0 23644 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1
transform -1 0 16376 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1
transform 1 0 48576 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1
transform -1 0 28796 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1
transform -1 0 13892 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1
transform -1 0 57224 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1
transform -1 0 40848 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1
transform -1 0 32844 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1
transform 1 0 30544 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1
transform 1 0 47012 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1
transform -1 0 46092 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1
transform -1 0 66148 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1
transform -1 0 60168 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1
transform -1 0 36616 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1
transform -1 0 36616 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1
transform -1 0 66148 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1
transform 1 0 47932 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1
transform 1 0 14628 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1
transform 1 0 59892 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1
transform -1 0 66148 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1
transform 1 0 48392 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1
transform -1 0 23736 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1
transform -1 0 57224 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1
transform -1 0 56396 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1
transform -1 0 41768 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1
transform -1 0 27968 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1
transform -1 0 35972 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1
transform -1 0 66148 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1
transform 1 0 47932 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1
transform 1 0 47104 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1
transform -1 0 41768 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1
transform -1 0 23644 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1
transform -1 0 12328 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1
transform -1 0 66148 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1
transform -1 0 65780 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1
transform 1 0 19228 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1
transform -1 0 40204 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1
transform -1 0 27140 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1
transform 1 0 34224 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1
transform 1 0 20424 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1
transform -1 0 9384 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1
transform 1 0 44896 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1
transform -1 0 43424 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1
transform -1 0 27968 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1
transform -1 0 30084 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1
transform -1 0 66148 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1
transform -1 0 52900 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1
transform -1 0 44620 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1
transform -1 0 20976 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1
transform -1 0 28612 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1
transform -1 0 11684 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1
transform -1 0 54280 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1
transform 1 0 10948 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1
transform -1 0 16008 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1
transform 1 0 43608 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1
transform -1 0 51980 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1
transform 1 0 18860 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1
transform -1 0 66148 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1
transform -1 0 16192 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1
transform -1 0 66148 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1
transform 1 0 38272 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1
transform -1 0 19412 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1
transform -1 0 34868 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1
transform -1 0 66148 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1
transform -1 0 18584 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1
transform -1 0 18768 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1
transform -1 0 40020 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1
transform -1 0 40020 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1
transform 1 0 31556 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1
transform -1 0 30544 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1
transform -1 0 28428 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1
transform -1 0 32384 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1
transform -1 0 34500 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1
transform -1 0 26220 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1
transform 1 0 23000 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1
transform 1 0 28612 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1
transform 1 0 26404 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1
transform -1 0 27508 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1
transform 1 0 26404 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_2_Left_66
timestamp 1
transform 1 0 63572 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_2_Right_147
timestamp 1
transform -1 0 66424 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_2_Left_0
timestamp 1
transform 1 0 63572 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_2_Right_67
timestamp 1
transform -1 0 66424 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_2_Left_1
timestamp 1
transform 1 0 63572 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_2_Right_68
timestamp 1
transform -1 0 66424 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_2_Left_2
timestamp 1
transform 1 0 63572 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_2_Right_69
timestamp 1
transform -1 0 66424 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_2_Left_3
timestamp 1
transform 1 0 63572 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_2_Right_70
timestamp 1
transform -1 0 66424 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_2_Left_4
timestamp 1
transform 1 0 63572 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_2_Right_71
timestamp 1
transform -1 0 66424 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_2_Left_5
timestamp 1
transform 1 0 63572 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_2_Right_72
timestamp 1
transform -1 0 66424 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_2_Left_6
timestamp 1
transform 1 0 63572 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_2_Right_73
timestamp 1
transform -1 0 66424 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_2_Left_7
timestamp 1
transform 1 0 63572 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_2_Right_74
timestamp 1
transform -1 0 66424 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_2_Left_8
timestamp 1
transform 1 0 63572 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_2_Right_75
timestamp 1
transform -1 0 66424 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Left_9
timestamp 1
transform 1 0 63572 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Right_76
timestamp 1
transform -1 0 66424 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Left_10
timestamp 1
transform 1 0 63572 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Right_77
timestamp 1
transform -1 0 66424 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Left_11
timestamp 1
transform 1 0 63572 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Right_78
timestamp 1
transform -1 0 66424 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Left_12
timestamp 1
transform 1 0 63572 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Right_79
timestamp 1
transform -1 0 66424 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Left_13
timestamp 1
transform 1 0 63572 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Right_80
timestamp 1
transform -1 0 66424 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Left_14
timestamp 1
transform 1 0 63572 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Right_81
timestamp 1
transform -1 0 66424 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Left_15
timestamp 1
transform 1 0 63572 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Right_82
timestamp 1
transform -1 0 66424 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Left_16
timestamp 1
transform 1 0 63572 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Right_83
timestamp 1
transform -1 0 66424 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Left_17
timestamp 1
transform 1 0 63572 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Right_84
timestamp 1
transform -1 0 66424 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Left_18
timestamp 1
transform 1 0 63572 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Right_85
timestamp 1
transform -1 0 66424 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Left_19
timestamp 1
transform 1 0 63572 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Right_86
timestamp 1
transform -1 0 66424 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Left_20
timestamp 1
transform 1 0 63572 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Right_87
timestamp 1
transform -1 0 66424 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Left_21
timestamp 1
transform 1 0 63572 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Right_88
timestamp 1
transform -1 0 66424 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Left_22
timestamp 1
transform 1 0 63572 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Right_89
timestamp 1
transform -1 0 66424 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Left_23
timestamp 1
transform 1 0 63572 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Right_90
timestamp 1
transform -1 0 66424 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Left_24
timestamp 1
transform 1 0 63572 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Right_91
timestamp 1
transform -1 0 66424 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Left_25
timestamp 1
transform 1 0 63572 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Right_92
timestamp 1
transform -1 0 66424 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Left_26
timestamp 1
transform 1 0 63572 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Right_93
timestamp 1
transform -1 0 66424 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Left_27
timestamp 1
transform 1 0 63572 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Right_94
timestamp 1
transform -1 0 66424 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Left_28
timestamp 1
transform 1 0 63572 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Right_95
timestamp 1
transform -1 0 66424 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Left_29
timestamp 1
transform 1 0 63572 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Right_96
timestamp 1
transform -1 0 66424 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Left_30
timestamp 1
transform 1 0 63572 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Right_97
timestamp 1
transform -1 0 66424 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Left_31
timestamp 1
transform 1 0 63572 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Right_98
timestamp 1
transform -1 0 66424 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Left_32
timestamp 1
transform 1 0 63572 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Right_99
timestamp 1
transform -1 0 66424 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Left_33
timestamp 1
transform 1 0 63572 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Right_100
timestamp 1
transform -1 0 66424 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Left_34
timestamp 1
transform 1 0 63572 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Right_101
timestamp 1
transform -1 0 66424 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Left_35
timestamp 1
transform 1 0 63572 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Right_102
timestamp 1
transform -1 0 66424 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Left_36
timestamp 1
transform 1 0 63572 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Right_103
timestamp 1
transform -1 0 66424 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Left_37
timestamp 1
transform 1 0 63572 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Right_104
timestamp 1
transform -1 0 66424 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Left_38
timestamp 1
transform 1 0 63572 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Right_105
timestamp 1
transform -1 0 66424 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Left_39
timestamp 1
transform 1 0 63572 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Right_106
timestamp 1
transform -1 0 66424 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Left_40
timestamp 1
transform 1 0 63572 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Right_107
timestamp 1
transform -1 0 66424 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Left_41
timestamp 1
transform 1 0 63572 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Right_108
timestamp 1
transform -1 0 66424 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Left_42
timestamp 1
transform 1 0 63572 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Right_109
timestamp 1
transform -1 0 66424 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Left_43
timestamp 1
transform 1 0 63572 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Right_110
timestamp 1
transform -1 0 66424 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Left_44
timestamp 1
transform 1 0 63572 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Right_111
timestamp 1
transform -1 0 66424 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Left_45
timestamp 1
transform 1 0 63572 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Right_112
timestamp 1
transform -1 0 66424 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Left_46
timestamp 1
transform 1 0 63572 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Right_113
timestamp 1
transform -1 0 66424 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Left_47
timestamp 1
transform 1 0 63572 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Right_114
timestamp 1
transform -1 0 66424 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Left_48
timestamp 1
transform 1 0 63572 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Right_115
timestamp 1
transform -1 0 66424 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Left_49
timestamp 1
transform 1 0 63572 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Right_116
timestamp 1
transform -1 0 66424 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Left_50
timestamp 1
transform 1 0 63572 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Right_117
timestamp 1
transform -1 0 66424 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Left_51
timestamp 1
transform 1 0 63572 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Right_118
timestamp 1
transform -1 0 66424 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Left_52
timestamp 1
transform 1 0 63572 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Right_119
timestamp 1
transform -1 0 66424 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Left_53
timestamp 1
transform 1 0 63572 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Right_120
timestamp 1
transform -1 0 66424 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Left_54
timestamp 1
transform 1 0 63572 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Right_121
timestamp 1
transform -1 0 66424 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Left_55
timestamp 1
transform 1 0 63572 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Right_122
timestamp 1
transform -1 0 66424 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Left_56
timestamp 1
transform 1 0 63572 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Right_123
timestamp 1
transform -1 0 66424 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Left_57
timestamp 1
transform 1 0 63572 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Right_124
timestamp 1
transform -1 0 66424 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Left_58
timestamp 1
transform 1 0 63572 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Right_125
timestamp 1
transform -1 0 66424 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Left_59
timestamp 1
transform 1 0 63572 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Right_126
timestamp 1
transform -1 0 66424 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Left_60
timestamp 1
transform 1 0 63572 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Right_127
timestamp 1
transform -1 0 66424 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Left_61
timestamp 1
transform 1 0 63572 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Right_128
timestamp 1
transform -1 0 66424 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Left_62
timestamp 1
transform 1 0 63572 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Right_129
timestamp 1
transform -1 0 66424 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Left_63
timestamp 1
transform 1 0 63572 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Right_130
timestamp 1
transform -1 0 66424 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Left_64
timestamp 1
transform 1 0 63572 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Right_131
timestamp 1
transform -1 0 66424 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Left_65
timestamp 1
transform 1 0 63572 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Right_132
timestamp 1
transform -1 0 66424 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_148
timestamp 1
transform 1 0 552 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_133
timestamp 1
transform -1 0 66424 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_149
timestamp 1
transform 1 0 552 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_134
timestamp 1
transform -1 0 66424 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Left_150
timestamp 1
transform 1 0 552 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Right_135
timestamp 1
transform -1 0 66424 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Left_151
timestamp 1
transform 1 0 552 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Right_136
timestamp 1
transform -1 0 66424 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Left_152
timestamp 1
transform 1 0 552 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Right_137
timestamp 1
transform -1 0 66424 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Left_153
timestamp 1
transform 1 0 552 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Right_138
timestamp 1
transform -1 0 66424 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Left_154
timestamp 1
transform 1 0 552 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Right_139
timestamp 1
transform -1 0 66424 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Left_155
timestamp 1
transform 1 0 552 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Right_140
timestamp 1
transform -1 0 66424 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Left_156
timestamp 1
transform 1 0 552 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Right_141
timestamp 1
transform -1 0 66424 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Left_157
timestamp 1
transform 1 0 552 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Right_142
timestamp 1
transform -1 0 66424 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Left_158
timestamp 1
transform 1 0 552 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Right_143
timestamp 1
transform -1 0 66424 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Left_159
timestamp 1
transform 1 0 552 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Right_144
timestamp 1
transform -1 0 66424 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Left_160
timestamp 1
transform 1 0 552 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Right_145
timestamp 1
transform -1 0 66424 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Left_161
timestamp 1
transform 1 0 552 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Right_146
timestamp 1
transform -1 0 66424 0 1 44064
box -38 -48 314 592
use sky130_sram_128B_1rw_32x32  SRAM
timestamp 0
transform -1 0 62536 0 -1 35514
box 0 0 1 1
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_162
timestamp 1
transform 1 0 3128 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_163
timestamp 1
transform 1 0 5704 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_164
timestamp 1
transform 1 0 8280 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_165
timestamp 1
transform 1 0 10856 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_166
timestamp 1
transform 1 0 13432 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_167
timestamp 1
transform 1 0 16008 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_168
timestamp 1
transform 1 0 18584 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_169
timestamp 1
transform 1 0 21160 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_170
timestamp 1
transform 1 0 23736 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_171
timestamp 1
transform 1 0 26312 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_172
timestamp 1
transform 1 0 28888 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_173
timestamp 1
transform 1 0 31464 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_174
timestamp 1
transform 1 0 34040 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_175
timestamp 1
transform 1 0 36616 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_176
timestamp 1
transform 1 0 39192 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_177
timestamp 1
transform 1 0 41768 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_178
timestamp 1
transform 1 0 44344 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_179
timestamp 1
transform 1 0 46920 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_180
timestamp 1
transform 1 0 49496 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_181
timestamp 1
transform 1 0 52072 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_182
timestamp 1
transform 1 0 54648 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_183
timestamp 1
transform 1 0 57224 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_184
timestamp 1
transform 1 0 59800 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_185
timestamp 1
transform 1 0 62376 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_186
timestamp 1
transform 1 0 64952 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_187
timestamp 1
transform 1 0 3128 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_188
timestamp 1
transform 1 0 8280 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_189
timestamp 1
transform 1 0 13432 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_190
timestamp 1
transform 1 0 18584 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_191
timestamp 1
transform 1 0 23736 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_192
timestamp 1
transform 1 0 28888 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_193
timestamp 1
transform 1 0 34040 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_194
timestamp 1
transform 1 0 39192 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_195
timestamp 1
transform 1 0 44344 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_196
timestamp 1
transform 1 0 49496 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_197
timestamp 1
transform 1 0 54648 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_198
timestamp 1
transform 1 0 59800 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_199
timestamp 1
transform 1 0 64952 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_200
timestamp 1
transform 1 0 5704 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_201
timestamp 1
transform 1 0 10856 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_202
timestamp 1
transform 1 0 16008 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_203
timestamp 1
transform 1 0 21160 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_204
timestamp 1
transform 1 0 26312 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_205
timestamp 1
transform 1 0 31464 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_206
timestamp 1
transform 1 0 36616 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_207
timestamp 1
transform 1 0 41768 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_208
timestamp 1
transform 1 0 46920 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_209
timestamp 1
transform 1 0 52072 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_210
timestamp 1
transform 1 0 57224 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_211
timestamp 1
transform 1 0 62376 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_212
timestamp 1
transform 1 0 3128 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_213
timestamp 1
transform 1 0 8280 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_214
timestamp 1
transform 1 0 13432 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_215
timestamp 1
transform 1 0 18584 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_216
timestamp 1
transform 1 0 23736 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_217
timestamp 1
transform 1 0 28888 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_218
timestamp 1
transform 1 0 34040 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_219
timestamp 1
transform 1 0 39192 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_220
timestamp 1
transform 1 0 44344 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_221
timestamp 1
transform 1 0 49496 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_222
timestamp 1
transform 1 0 54648 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_223
timestamp 1
transform 1 0 59800 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_224
timestamp 1
transform 1 0 64952 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_225
timestamp 1
transform 1 0 5704 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_226
timestamp 1
transform 1 0 10856 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_227
timestamp 1
transform 1 0 16008 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_228
timestamp 1
transform 1 0 21160 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_229
timestamp 1
transform 1 0 26312 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_230
timestamp 1
transform 1 0 31464 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_231
timestamp 1
transform 1 0 36616 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_232
timestamp 1
transform 1 0 41768 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_233
timestamp 1
transform 1 0 46920 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_234
timestamp 1
transform 1 0 52072 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_235
timestamp 1
transform 1 0 57224 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_236
timestamp 1
transform 1 0 62376 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_237
timestamp 1
transform 1 0 3128 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_238
timestamp 1
transform 1 0 8280 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_239
timestamp 1
transform 1 0 13432 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_240
timestamp 1
transform 1 0 18584 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_241
timestamp 1
transform 1 0 23736 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_242
timestamp 1
transform 1 0 28888 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_243
timestamp 1
transform 1 0 34040 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_244
timestamp 1
transform 1 0 39192 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_245
timestamp 1
transform 1 0 44344 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_246
timestamp 1
transform 1 0 49496 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_247
timestamp 1
transform 1 0 54648 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_248
timestamp 1
transform 1 0 59800 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_249
timestamp 1
transform 1 0 64952 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_250
timestamp 1
transform 1 0 5704 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_251
timestamp 1
transform 1 0 10856 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_252
timestamp 1
transform 1 0 16008 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_253
timestamp 1
transform 1 0 21160 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_254
timestamp 1
transform 1 0 26312 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_255
timestamp 1
transform 1 0 31464 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_256
timestamp 1
transform 1 0 36616 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_257
timestamp 1
transform 1 0 41768 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_258
timestamp 1
transform 1 0 46920 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_259
timestamp 1
transform 1 0 52072 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_260
timestamp 1
transform 1 0 57224 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_261
timestamp 1
transform 1 0 62376 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_262
timestamp 1
transform 1 0 3128 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_263
timestamp 1
transform 1 0 8280 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_264
timestamp 1
transform 1 0 13432 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_265
timestamp 1
transform 1 0 18584 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_266
timestamp 1
transform 1 0 23736 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_267
timestamp 1
transform 1 0 28888 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_268
timestamp 1
transform 1 0 34040 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_269
timestamp 1
transform 1 0 39192 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_270
timestamp 1
transform 1 0 44344 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_271
timestamp 1
transform 1 0 49496 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_272
timestamp 1
transform 1 0 54648 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_273
timestamp 1
transform 1 0 59800 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_274
timestamp 1
transform 1 0 64952 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_275
timestamp 1
transform 1 0 5704 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_276
timestamp 1
transform 1 0 10856 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_277
timestamp 1
transform 1 0 16008 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_278
timestamp 1
transform 1 0 21160 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_279
timestamp 1
transform 1 0 26312 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_280
timestamp 1
transform 1 0 31464 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_281
timestamp 1
transform 1 0 36616 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_282
timestamp 1
transform 1 0 41768 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_283
timestamp 1
transform 1 0 46920 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_284
timestamp 1
transform 1 0 52072 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_285
timestamp 1
transform 1 0 57224 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_286
timestamp 1
transform 1 0 62376 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_287
timestamp 1
transform 1 0 3128 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_288
timestamp 1
transform 1 0 8280 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_289
timestamp 1
transform 1 0 13432 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_290
timestamp 1
transform 1 0 18584 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_291
timestamp 1
transform 1 0 23736 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_292
timestamp 1
transform 1 0 28888 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_293
timestamp 1
transform 1 0 34040 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_294
timestamp 1
transform 1 0 39192 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_295
timestamp 1
transform 1 0 44344 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_296
timestamp 1
transform 1 0 49496 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_297
timestamp 1
transform 1 0 54648 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_298
timestamp 1
transform 1 0 59800 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_299
timestamp 1
transform 1 0 64952 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_300
timestamp 1
transform 1 0 5704 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_301
timestamp 1
transform 1 0 10856 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_302
timestamp 1
transform 1 0 16008 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_303
timestamp 1
transform 1 0 21160 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_304
timestamp 1
transform 1 0 26312 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_305
timestamp 1
transform 1 0 31464 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_306
timestamp 1
transform 1 0 36616 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_307
timestamp 1
transform 1 0 41768 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_308
timestamp 1
transform 1 0 46920 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_309
timestamp 1
transform 1 0 52072 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_310
timestamp 1
transform 1 0 57224 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_311
timestamp 1
transform 1 0 62376 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_312
timestamp 1
transform 1 0 3128 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_313
timestamp 1
transform 1 0 8280 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_314
timestamp 1
transform 1 0 13432 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_315
timestamp 1
transform 1 0 18584 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_316
timestamp 1
transform 1 0 23736 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_317
timestamp 1
transform 1 0 28888 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_318
timestamp 1
transform 1 0 34040 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_319
timestamp 1
transform 1 0 39192 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_320
timestamp 1
transform 1 0 44344 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_321
timestamp 1
transform 1 0 49496 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_322
timestamp 1
transform 1 0 54648 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_323
timestamp 1
transform 1 0 59800 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_324
timestamp 1
transform 1 0 64952 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_325
timestamp 1
transform 1 0 5704 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_326
timestamp 1
transform 1 0 10856 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_327
timestamp 1
transform 1 0 16008 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_328
timestamp 1
transform 1 0 21160 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_329
timestamp 1
transform 1 0 26312 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_330
timestamp 1
transform 1 0 31464 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_331
timestamp 1
transform 1 0 36616 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_332
timestamp 1
transform 1 0 41768 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_333
timestamp 1
transform 1 0 46920 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_334
timestamp 1
transform 1 0 52072 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_335
timestamp 1
transform 1 0 57224 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_336
timestamp 1
transform 1 0 62376 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_337
timestamp 1
transform 1 0 3128 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_338
timestamp 1
transform 1 0 5704 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_339
timestamp 1
transform 1 0 8280 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_340
timestamp 1
transform 1 0 10856 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_341
timestamp 1
transform 1 0 13432 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_342
timestamp 1
transform 1 0 16008 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_343
timestamp 1
transform 1 0 18584 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_344
timestamp 1
transform 1 0 21160 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_345
timestamp 1
transform 1 0 23736 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_346
timestamp 1
transform 1 0 26312 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_347
timestamp 1
transform 1 0 28888 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_348
timestamp 1
transform 1 0 31464 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_349
timestamp 1
transform 1 0 34040 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_350
timestamp 1
transform 1 0 36616 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_351
timestamp 1
transform 1 0 39192 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_352
timestamp 1
transform 1 0 41768 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_353
timestamp 1
transform 1 0 44344 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_354
timestamp 1
transform 1 0 46920 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_355
timestamp 1
transform 1 0 49496 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_356
timestamp 1
transform 1 0 52072 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_357
timestamp 1
transform 1 0 54648 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_358
timestamp 1
transform 1 0 57224 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_359
timestamp 1
transform 1 0 59800 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_360
timestamp 1
transform 1 0 62376 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_361
timestamp 1
transform 1 0 64952 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_56
timestamp 1
transform -1 0 10304 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_57
timestamp 1
transform -1 0 9752 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_58
timestamp 1
transform -1 0 9200 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_59
timestamp 1
transform -1 0 8648 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_60
timestamp 1
transform -1 0 8096 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_61
timestamp 1
transform -1 0 7544 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_62
timestamp 1
transform -1 0 6992 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_63
timestamp 1
transform -1 0 6440 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_64
timestamp 1
transform -1 0 15548 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_65
timestamp 1
transform -1 0 14076 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_66
timestamp 1
transform -1 0 13800 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_67
timestamp 1
transform -1 0 13064 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_68
timestamp 1
transform -1 0 12512 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_69
timestamp 1
transform -1 0 12788 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_70
timestamp 1
transform -1 0 11408 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_71
timestamp 1
transform -1 0 10856 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_72
timestamp 1
transform 1 0 17020 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_73
timestamp 1
transform 1 0 16744 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_74
timestamp 1
transform 1 0 16468 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_75
timestamp 1
transform 1 0 15732 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_76
timestamp 1
transform -1 0 15732 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_openram_top_77
timestamp 1
transform -1 0 16468 0 1 44064
box -38 -48 314 592
<< labels >>
flabel metal4 s 2912 34210 3232 44656 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 51912 34142 52232 44656 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 65252 496 65572 37584 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1992 34208 2312 44656 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 50992 34142 51312 44656 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 64332 496 64652 37584 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 2 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 3 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 4 nsew signal input
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 5 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 6 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 7 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 8 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 9 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 10 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 11 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 12 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 13 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 14 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 15 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 16 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 17 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 18 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 19 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 20 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 21 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 22 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 23 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 24 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 25 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 26 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 27 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 28 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 29 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 30 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 31 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 32 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 33 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 34 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 35 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 36 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 37 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 38 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 39 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 40 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 41 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 42 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 43 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 44 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 66976 45152
<< end >>
