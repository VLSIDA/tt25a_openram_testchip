module tt_um_openram_top (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire \dout[0] ;
 wire \dout[10] ;
 wire \dout[11] ;
 wire \dout[12] ;
 wire \dout[13] ;
 wire \dout[14] ;
 wire \dout[15] ;
 wire \dout[16] ;
 wire \dout[17] ;
 wire \dout[18] ;
 wire \dout[19] ;
 wire \dout[1] ;
 wire \dout[20] ;
 wire \dout[21] ;
 wire \dout[22] ;
 wire \dout[23] ;
 wire \dout[24] ;
 wire \dout[25] ;
 wire \dout[26] ;
 wire \dout[27] ;
 wire \dout[28] ;
 wire \dout[29] ;
 wire \dout[2] ;
 wire \dout[30] ;
 wire \dout[31] ;
 wire \dout[32] ;
 wire \dout[3] ;
 wire \dout[4] ;
 wire \dout[5] ;
 wire \dout[6] ;
 wire \dout[7] ;
 wire \dout[8] ;
 wire \dout[9] ;
 wire \scan_chain.scan_cells[0].scan_cell.data_out ;
 wire \scan_chain.scan_cells[0].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[10].scan_cell.data_out ;
 wire \scan_chain.scan_cells[10].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[10].scan_cell.scan_in ;
 wire \scan_chain.scan_cells[11].scan_cell.data_out ;
 wire \scan_chain.scan_cells[11].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[12].scan_cell.data_out ;
 wire \scan_chain.scan_cells[12].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[13].scan_cell.data_out ;
 wire \scan_chain.scan_cells[13].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[14].scan_cell.data_out ;
 wire \scan_chain.scan_cells[14].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[15].scan_cell.data_out ;
 wire \scan_chain.scan_cells[15].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[16].scan_cell.data_out ;
 wire \scan_chain.scan_cells[16].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[17].scan_cell.data_out ;
 wire \scan_chain.scan_cells[17].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[18].scan_cell.data_out ;
 wire \scan_chain.scan_cells[18].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[19].scan_cell.data_out ;
 wire \scan_chain.scan_cells[19].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[1].scan_cell.data_out ;
 wire \scan_chain.scan_cells[1].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[20].scan_cell.data_out ;
 wire \scan_chain.scan_cells[20].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[21].scan_cell.data_out ;
 wire \scan_chain.scan_cells[21].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[22].scan_cell.data_out ;
 wire \scan_chain.scan_cells[22].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[23].scan_cell.data_out ;
 wire \scan_chain.scan_cells[23].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[24].scan_cell.data_out ;
 wire \scan_chain.scan_cells[24].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[25].scan_cell.data_out ;
 wire \scan_chain.scan_cells[25].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[26].scan_cell.data_out ;
 wire \scan_chain.scan_cells[26].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[27].scan_cell.data_out ;
 wire \scan_chain.scan_cells[27].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[28].scan_cell.data_out ;
 wire \scan_chain.scan_cells[28].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[29].scan_cell.data_out ;
 wire \scan_chain.scan_cells[29].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[2].scan_cell.data_out ;
 wire \scan_chain.scan_cells[2].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[30].scan_cell.data_out ;
 wire \scan_chain.scan_cells[30].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[31].scan_cell.data_out ;
 wire \scan_chain.scan_cells[31].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[32].scan_cell.data_out ;
 wire \scan_chain.scan_cells[32].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[33].scan_cell.data_in ;
 wire \scan_chain.scan_cells[33].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[34].scan_cell.data_in ;
 wire \scan_chain.scan_cells[34].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[35].scan_cell.data_in ;
 wire \scan_chain.scan_cells[35].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[36].scan_cell.data_in ;
 wire \scan_chain.scan_cells[36].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[37].scan_cell.data_in ;
 wire \scan_chain.scan_cells[37].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[38].scan_cell.data_in ;
 wire \scan_chain.scan_cells[38].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[39].scan_cell.data_in ;
 wire \scan_chain.scan_cells[39].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[3].scan_cell.data_out ;
 wire \scan_chain.scan_cells[3].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[40].scan_cell.data_in ;
 wire \scan_chain.scan_cells[40].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[41].scan_cell.data_in ;
 wire \scan_chain.scan_cells[41].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[42].scan_cell.data_in ;
 wire \scan_chain.scan_cells[42].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[43].scan_cell.data_in ;
 wire \scan_chain.scan_cells[43].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[44].scan_cell.data_in ;
 wire \scan_chain.scan_cells[44].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[45].scan_cell.data_in ;
 wire \scan_chain.scan_cells[45].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[46].scan_cell.data_in ;
 wire \scan_chain.scan_cells[46].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[47].scan_cell.data_in ;
 wire \scan_chain.scan_cells[47].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[48].scan_cell.data_in ;
 wire \scan_chain.scan_cells[48].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[49].scan_cell.data_in ;
 wire \scan_chain.scan_cells[49].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[4].scan_cell.data_out ;
 wire \scan_chain.scan_cells[4].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[50].scan_cell.data_in ;
 wire \scan_chain.scan_cells[50].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[51].scan_cell.data_in ;
 wire \scan_chain.scan_cells[51].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[52].scan_cell.data_in ;
 wire \scan_chain.scan_cells[52].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[53].scan_cell.data_in ;
 wire \scan_chain.scan_cells[53].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[54].scan_cell.data_in ;
 wire \scan_chain.scan_cells[54].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[55].scan_cell.data_in ;
 wire \scan_chain.scan_cells[55].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[56].scan_cell.data_in ;
 wire \scan_chain.scan_cells[56].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[57].scan_cell.data_in ;
 wire \scan_chain.scan_cells[57].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[58].scan_cell.data_in ;
 wire \scan_chain.scan_cells[58].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[59].scan_cell.data_in ;
 wire \scan_chain.scan_cells[59].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[5].scan_cell.data_out ;
 wire \scan_chain.scan_cells[5].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[60].scan_cell.data_in ;
 wire \scan_chain.scan_cells[60].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[61].scan_cell.data_in ;
 wire \scan_chain.scan_cells[61].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[62].scan_cell.data_in ;
 wire \scan_chain.scan_cells[62].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[63].scan_cell.data_in ;
 wire \scan_chain.scan_cells[63].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[64].scan_cell.data_in ;
 wire \scan_chain.scan_cells[64].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[65].scan_cell.data_in ;
 wire \scan_chain.scan_cells[65].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[66].scan_cell.data_in ;
 wire \scan_chain.scan_cells[66].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[67].scan_cell.data_in ;
 wire \scan_chain.scan_cells[67].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[68].scan_cell.data_in ;
 wire \scan_chain.scan_cells[68].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[69].scan_cell.data_in ;
 wire \scan_chain.scan_cells[69].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[6].scan_cell.data_out ;
 wire \scan_chain.scan_cells[6].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[70].scan_cell.data_in ;
 wire \scan_chain.scan_cells[70].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[71].scan_cell.data_in ;
 wire \scan_chain.scan_cells[71].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[7].scan_cell.data_out ;
 wire \scan_chain.scan_cells[7].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[8].scan_cell.data_out ;
 wire \scan_chain.scan_cells[8].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[9].scan_cell.primary_ff ;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire vccd1;
 wire vssd1;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire [4:0] clknet_0_ui_in;
 wire [4:0] clknet_3_0__leaf_ui_in;
 wire [4:0] clknet_3_1__leaf_ui_in;
 wire [4:0] clknet_3_2__leaf_ui_in;
 wire [4:0] clknet_3_3__leaf_ui_in;
 wire [4:0] clknet_3_4__leaf_ui_in;
 wire [4:0] clknet_3_5__leaf_ui_in;
 wire [4:0] clknet_3_6__leaf_ui_in;
 wire [4:0] clknet_3_7__leaf_ui_in;

 sky130_sram_128B_1rw_32x32 SRAM (.csb0(ui_in[5]),
    .web0(ui_in[6]),
    .clk0(clknet_3_4__leaf_ui_in[3]),
    .spare_wen0(ui_in[7]),
    .vccd1(VPWR),
    .vssd1(VGND),
    .addr0({\scan_chain.scan_cells[71].scan_cell.data_in ,
    \scan_chain.scan_cells[70].scan_cell.data_in ,
    \scan_chain.scan_cells[69].scan_cell.data_in ,
    \scan_chain.scan_cells[68].scan_cell.data_in ,
    \scan_chain.scan_cells[67].scan_cell.data_in ,
    \scan_chain.scan_cells[66].scan_cell.data_in }),
    .din0({\scan_chain.scan_cells[65].scan_cell.data_in ,
    \scan_chain.scan_cells[64].scan_cell.data_in ,
    \scan_chain.scan_cells[63].scan_cell.data_in ,
    \scan_chain.scan_cells[62].scan_cell.data_in ,
    \scan_chain.scan_cells[61].scan_cell.data_in ,
    \scan_chain.scan_cells[60].scan_cell.data_in ,
    \scan_chain.scan_cells[59].scan_cell.data_in ,
    \scan_chain.scan_cells[58].scan_cell.data_in ,
    \scan_chain.scan_cells[57].scan_cell.data_in ,
    \scan_chain.scan_cells[56].scan_cell.data_in ,
    \scan_chain.scan_cells[55].scan_cell.data_in ,
    \scan_chain.scan_cells[54].scan_cell.data_in ,
    \scan_chain.scan_cells[53].scan_cell.data_in ,
    \scan_chain.scan_cells[52].scan_cell.data_in ,
    \scan_chain.scan_cells[51].scan_cell.data_in ,
    \scan_chain.scan_cells[50].scan_cell.data_in ,
    \scan_chain.scan_cells[49].scan_cell.data_in ,
    \scan_chain.scan_cells[48].scan_cell.data_in ,
    \scan_chain.scan_cells[47].scan_cell.data_in ,
    \scan_chain.scan_cells[46].scan_cell.data_in ,
    \scan_chain.scan_cells[45].scan_cell.data_in ,
    \scan_chain.scan_cells[44].scan_cell.data_in ,
    \scan_chain.scan_cells[43].scan_cell.data_in ,
    \scan_chain.scan_cells[42].scan_cell.data_in ,
    \scan_chain.scan_cells[41].scan_cell.data_in ,
    \scan_chain.scan_cells[40].scan_cell.data_in ,
    \scan_chain.scan_cells[39].scan_cell.data_in ,
    \scan_chain.scan_cells[38].scan_cell.data_in ,
    \scan_chain.scan_cells[37].scan_cell.data_in ,
    \scan_chain.scan_cells[36].scan_cell.data_in ,
    \scan_chain.scan_cells[35].scan_cell.data_in ,
    \scan_chain.scan_cells[34].scan_cell.data_in ,
    \scan_chain.scan_cells[33].scan_cell.data_in }),
    .dout0({\dout[32] ,
    \dout[31] ,
    \dout[30] ,
    \dout[29] ,
    \dout[28] ,
    \dout[27] ,
    \dout[26] ,
    \dout[25] ,
    \dout[24] ,
    \dout[23] ,
    \dout[22] ,
    \dout[21] ,
    \dout[20] ,
    \dout[19] ,
    \dout[18] ,
    \dout[17] ,
    \dout[16] ,
    \dout[15] ,
    \dout[14] ,
    \dout[13] ,
    \dout[12] ,
    \dout[11] ,
    \dout[10] ,
    \dout[9] ,
    \dout[8] ,
    \dout[7] ,
    \dout[6] ,
    \dout[5] ,
    \dout[4] ,
    \dout[3] ,
    \dout[2] ,
    \dout[1] ,
    \dout[0] }),
    .wmask0({uio_in[3],
    uio_in[2],
    uio_in[1],
    uio_in[0]}));
 sky130_fd_sc_hd__mux2_1 _250_ (.A0(\scan_chain.scan_cells[10].scan_cell.scan_in ),
    .A1(\scan_chain.scan_cells[8].scan_cell.data_out ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_144_));
 sky130_fd_sc_hd__mux2_1 _251_ (.A0(\scan_chain.scan_cells[9].scan_cell.primary_ff ),
    .A1(_144_),
    .S(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_026_));
 sky130_fd_sc_hd__nand2_2 _252_ (.A(net21),
    .B(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_145_));
 sky130_fd_sc_hd__mux2_1 _253_ (.A0(\scan_chain.scan_cells[71].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[71].scan_cell.data_in ),
    .S(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_027_));
 sky130_fd_sc_hd__mux2_1 _254_ (.A0(\scan_chain.scan_cells[70].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[69].scan_cell.data_in ),
    .S(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_146_));
 sky130_fd_sc_hd__mux2_1 _255_ (.A0(\scan_chain.scan_cells[70].scan_cell.primary_ff ),
    .A1(_146_),
    .S(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_028_));
 sky130_fd_sc_hd__mux2_1 _256_ (.A0(\scan_chain.scan_cells[70].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[70].scan_cell.data_in ),
    .S(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _257_ (.A0(\scan_chain.scan_cells[6].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[5].scan_cell.data_out ),
    .S(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_147_));
 sky130_fd_sc_hd__mux2_1 _258_ (.A0(\scan_chain.scan_cells[6].scan_cell.primary_ff ),
    .A1(_147_),
    .S(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _259_ (.A0(\scan_chain.scan_cells[69].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[69].scan_cell.data_in ),
    .S(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_031_));
 sky130_fd_sc_hd__mux2_1 _260_ (.A0(\scan_chain.scan_cells[68].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[67].scan_cell.data_in ),
    .S(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_148_));
 sky130_fd_sc_hd__mux2_1 _261_ (.A0(\scan_chain.scan_cells[68].scan_cell.primary_ff ),
    .A1(_148_),
    .S(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_032_));
 sky130_fd_sc_hd__mux2_1 _262_ (.A0(\scan_chain.scan_cells[68].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[68].scan_cell.data_in ),
    .S(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_033_));
 sky130_fd_sc_hd__mux2_1 _263_ (.A0(\scan_chain.scan_cells[67].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[66].scan_cell.data_in ),
    .S(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_149_));
 sky130_fd_sc_hd__mux2_1 _264_ (.A0(\scan_chain.scan_cells[67].scan_cell.primary_ff ),
    .A1(_149_),
    .S(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_034_));
 sky130_fd_sc_hd__mux2_1 _265_ (.A0(\scan_chain.scan_cells[67].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[67].scan_cell.data_in ),
    .S(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_035_));
 sky130_fd_sc_hd__mux2_1 _266_ (.A0(\scan_chain.scan_cells[66].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[65].scan_cell.data_in ),
    .S(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_150_));
 sky130_fd_sc_hd__mux2_1 _267_ (.A0(\scan_chain.scan_cells[66].scan_cell.primary_ff ),
    .A1(_150_),
    .S(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_036_));
 sky130_fd_sc_hd__mux2_1 _268_ (.A0(\scan_chain.scan_cells[66].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[66].scan_cell.data_in ),
    .S(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_037_));
 sky130_fd_sc_hd__mux2_1 _269_ (.A0(\scan_chain.scan_cells[65].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[64].scan_cell.data_in ),
    .S(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_151_));
 sky130_fd_sc_hd__mux2_1 _270_ (.A0(\scan_chain.scan_cells[65].scan_cell.primary_ff ),
    .A1(_151_),
    .S(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_038_));
 sky130_fd_sc_hd__mux2_1 _271_ (.A0(\scan_chain.scan_cells[65].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[65].scan_cell.data_in ),
    .S(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_039_));
 sky130_fd_sc_hd__mux2_1 _272_ (.A0(\scan_chain.scan_cells[64].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[63].scan_cell.data_in ),
    .S(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_152_));
 sky130_fd_sc_hd__mux2_1 _273_ (.A0(\scan_chain.scan_cells[64].scan_cell.primary_ff ),
    .A1(_152_),
    .S(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_040_));
 sky130_fd_sc_hd__mux2_1 _274_ (.A0(\scan_chain.scan_cells[64].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[64].scan_cell.data_in ),
    .S(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_041_));
 sky130_fd_sc_hd__mux2_1 _275_ (.A0(\scan_chain.scan_cells[63].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[62].scan_cell.data_in ),
    .S(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_153_));
 sky130_fd_sc_hd__mux2_1 _276_ (.A0(\scan_chain.scan_cells[63].scan_cell.primary_ff ),
    .A1(_153_),
    .S(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_042_));
 sky130_fd_sc_hd__mux2_1 _277_ (.A0(\scan_chain.scan_cells[63].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[63].scan_cell.data_in ),
    .S(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_043_));
 sky130_fd_sc_hd__mux2_1 _278_ (.A0(\scan_chain.scan_cells[62].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[61].scan_cell.data_in ),
    .S(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_154_));
 sky130_fd_sc_hd__mux2_1 _279_ (.A0(\scan_chain.scan_cells[62].scan_cell.primary_ff ),
    .A1(_154_),
    .S(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_044_));
 sky130_fd_sc_hd__mux2_1 _280_ (.A0(\scan_chain.scan_cells[62].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[62].scan_cell.data_in ),
    .S(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_045_));
 sky130_fd_sc_hd__mux2_1 _281_ (.A0(\scan_chain.scan_cells[61].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[60].scan_cell.data_in ),
    .S(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_155_));
 sky130_fd_sc_hd__mux2_1 _282_ (.A0(\scan_chain.scan_cells[61].scan_cell.primary_ff ),
    .A1(_155_),
    .S(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_046_));
 sky130_fd_sc_hd__mux2_1 _283_ (.A0(\scan_chain.scan_cells[61].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[61].scan_cell.data_in ),
    .S(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_047_));
 sky130_fd_sc_hd__mux2_1 _284_ (.A0(\scan_chain.scan_cells[60].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[59].scan_cell.data_in ),
    .S(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_156_));
 sky130_fd_sc_hd__mux2_1 _285_ (.A0(\scan_chain.scan_cells[60].scan_cell.primary_ff ),
    .A1(_156_),
    .S(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_048_));
 sky130_fd_sc_hd__mux2_1 _286_ (.A0(\scan_chain.scan_cells[60].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[60].scan_cell.data_in ),
    .S(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_049_));
 sky130_fd_sc_hd__mux2_1 _287_ (.A0(\scan_chain.scan_cells[5].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[4].scan_cell.data_out ),
    .S(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_157_));
 sky130_fd_sc_hd__mux2_1 _288_ (.A0(\scan_chain.scan_cells[5].scan_cell.primary_ff ),
    .A1(_157_),
    .S(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_050_));
 sky130_fd_sc_hd__mux2_1 _289_ (.A0(\scan_chain.scan_cells[59].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[59].scan_cell.data_in ),
    .S(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_051_));
 sky130_fd_sc_hd__mux2_1 _290_ (.A0(\scan_chain.scan_cells[58].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[57].scan_cell.data_in ),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_158_));
 sky130_fd_sc_hd__mux2_1 _291_ (.A0(\scan_chain.scan_cells[58].scan_cell.primary_ff ),
    .A1(_158_),
    .S(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_052_));
 sky130_fd_sc_hd__mux2_1 _292_ (.A0(\scan_chain.scan_cells[58].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[58].scan_cell.data_in ),
    .S(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_053_));
 sky130_fd_sc_hd__mux2_1 _293_ (.A0(\scan_chain.scan_cells[57].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[56].scan_cell.data_in ),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_159_));
 sky130_fd_sc_hd__mux2_1 _294_ (.A0(\scan_chain.scan_cells[57].scan_cell.primary_ff ),
    .A1(_159_),
    .S(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_054_));
 sky130_fd_sc_hd__mux2_1 _295_ (.A0(\scan_chain.scan_cells[57].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[57].scan_cell.data_in ),
    .S(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_055_));
 sky130_fd_sc_hd__mux2_1 _296_ (.A0(\scan_chain.scan_cells[56].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[55].scan_cell.data_in ),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_160_));
 sky130_fd_sc_hd__mux2_1 _297_ (.A0(\scan_chain.scan_cells[56].scan_cell.primary_ff ),
    .A1(_160_),
    .S(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_056_));
 sky130_fd_sc_hd__mux2_1 _298_ (.A0(\scan_chain.scan_cells[56].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[56].scan_cell.data_in ),
    .S(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_057_));
 sky130_fd_sc_hd__mux2_1 _299_ (.A0(\scan_chain.scan_cells[55].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[54].scan_cell.data_in ),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_161_));
 sky130_fd_sc_hd__mux2_1 _300_ (.A0(\scan_chain.scan_cells[55].scan_cell.primary_ff ),
    .A1(_161_),
    .S(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_058_));
 sky130_fd_sc_hd__mux2_1 _301_ (.A0(\scan_chain.scan_cells[55].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[55].scan_cell.data_in ),
    .S(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_059_));
 sky130_fd_sc_hd__mux2_1 _302_ (.A0(\scan_chain.scan_cells[54].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[53].scan_cell.data_in ),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_162_));
 sky130_fd_sc_hd__mux2_1 _303_ (.A0(\scan_chain.scan_cells[54].scan_cell.primary_ff ),
    .A1(_162_),
    .S(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_060_));
 sky130_fd_sc_hd__mux2_1 _304_ (.A0(\scan_chain.scan_cells[54].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[54].scan_cell.data_in ),
    .S(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_061_));
 sky130_fd_sc_hd__mux2_1 _305_ (.A0(\scan_chain.scan_cells[53].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[52].scan_cell.data_in ),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_163_));
 sky130_fd_sc_hd__mux2_1 _306_ (.A0(\scan_chain.scan_cells[53].scan_cell.primary_ff ),
    .A1(_163_),
    .S(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_062_));
 sky130_fd_sc_hd__mux2_1 _307_ (.A0(\scan_chain.scan_cells[53].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[53].scan_cell.data_in ),
    .S(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_063_));
 sky130_fd_sc_hd__mux2_1 _308_ (.A0(\scan_chain.scan_cells[52].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[51].scan_cell.data_in ),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_164_));
 sky130_fd_sc_hd__mux2_1 _309_ (.A0(\scan_chain.scan_cells[52].scan_cell.primary_ff ),
    .A1(_164_),
    .S(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_064_));
 sky130_fd_sc_hd__mux2_1 _310_ (.A0(\scan_chain.scan_cells[52].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[52].scan_cell.data_in ),
    .S(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_065_));
 sky130_fd_sc_hd__mux2_1 _311_ (.A0(\scan_chain.scan_cells[51].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[50].scan_cell.data_in ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_165_));
 sky130_fd_sc_hd__mux2_1 _312_ (.A0(\scan_chain.scan_cells[51].scan_cell.primary_ff ),
    .A1(_165_),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_066_));
 sky130_fd_sc_hd__mux2_1 _313_ (.A0(\scan_chain.scan_cells[51].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[51].scan_cell.data_in ),
    .S(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_067_));
 sky130_fd_sc_hd__mux2_1 _314_ (.A0(\scan_chain.scan_cells[50].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[49].scan_cell.data_in ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_166_));
 sky130_fd_sc_hd__mux2_1 _315_ (.A0(\scan_chain.scan_cells[50].scan_cell.primary_ff ),
    .A1(_166_),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_068_));
 sky130_fd_sc_hd__mux2_1 _316_ (.A0(\scan_chain.scan_cells[50].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[50].scan_cell.data_in ),
    .S(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_069_));
 sky130_fd_sc_hd__mux2_1 _317_ (.A0(\scan_chain.scan_cells[4].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[3].scan_cell.data_out ),
    .S(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_167_));
 sky130_fd_sc_hd__mux2_1 _318_ (.A0(\scan_chain.scan_cells[4].scan_cell.primary_ff ),
    .A1(_167_),
    .S(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_070_));
 sky130_fd_sc_hd__mux2_1 _319_ (.A0(\scan_chain.scan_cells[49].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[49].scan_cell.data_in ),
    .S(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_071_));
 sky130_fd_sc_hd__mux2_1 _320_ (.A0(\scan_chain.scan_cells[48].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[47].scan_cell.data_in ),
    .S(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_168_));
 sky130_fd_sc_hd__mux2_1 _321_ (.A0(\scan_chain.scan_cells[48].scan_cell.primary_ff ),
    .A1(_168_),
    .S(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_072_));
 sky130_fd_sc_hd__mux2_1 _322_ (.A0(\scan_chain.scan_cells[48].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[48].scan_cell.data_in ),
    .S(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_073_));
 sky130_fd_sc_hd__mux2_1 _323_ (.A0(\scan_chain.scan_cells[47].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[46].scan_cell.data_in ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_169_));
 sky130_fd_sc_hd__mux2_1 _324_ (.A0(\scan_chain.scan_cells[47].scan_cell.primary_ff ),
    .A1(_169_),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_074_));
 sky130_fd_sc_hd__mux2_1 _325_ (.A0(\scan_chain.scan_cells[47].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[47].scan_cell.data_in ),
    .S(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_075_));
 sky130_fd_sc_hd__mux2_1 _326_ (.A0(\scan_chain.scan_cells[46].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[45].scan_cell.data_in ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_170_));
 sky130_fd_sc_hd__mux2_1 _327_ (.A0(\scan_chain.scan_cells[46].scan_cell.primary_ff ),
    .A1(_170_),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_076_));
 sky130_fd_sc_hd__mux2_1 _328_ (.A0(\scan_chain.scan_cells[46].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[46].scan_cell.data_in ),
    .S(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_077_));
 sky130_fd_sc_hd__mux2_1 _329_ (.A0(\scan_chain.scan_cells[45].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[44].scan_cell.data_in ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_171_));
 sky130_fd_sc_hd__mux2_1 _330_ (.A0(\scan_chain.scan_cells[45].scan_cell.primary_ff ),
    .A1(_171_),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_078_));
 sky130_fd_sc_hd__mux2_1 _331_ (.A0(\scan_chain.scan_cells[45].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[45].scan_cell.data_in ),
    .S(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_079_));
 sky130_fd_sc_hd__mux2_1 _332_ (.A0(\scan_chain.scan_cells[44].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[43].scan_cell.data_in ),
    .S(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_172_));
 sky130_fd_sc_hd__mux2_1 _333_ (.A0(\scan_chain.scan_cells[44].scan_cell.primary_ff ),
    .A1(_172_),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_080_));
 sky130_fd_sc_hd__mux2_1 _334_ (.A0(\scan_chain.scan_cells[44].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[44].scan_cell.data_in ),
    .S(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_081_));
 sky130_fd_sc_hd__mux2_1 _335_ (.A0(\scan_chain.scan_cells[43].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[42].scan_cell.data_in ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_173_));
 sky130_fd_sc_hd__mux2_1 _336_ (.A0(\scan_chain.scan_cells[43].scan_cell.primary_ff ),
    .A1(_173_),
    .S(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_082_));
 sky130_fd_sc_hd__mux2_1 _337_ (.A0(\scan_chain.scan_cells[43].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[43].scan_cell.data_in ),
    .S(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_083_));
 sky130_fd_sc_hd__mux2_1 _338_ (.A0(\scan_chain.scan_cells[42].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[41].scan_cell.data_in ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_174_));
 sky130_fd_sc_hd__mux2_1 _339_ (.A0(\scan_chain.scan_cells[42].scan_cell.primary_ff ),
    .A1(_174_),
    .S(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_084_));
 sky130_fd_sc_hd__mux2_1 _340_ (.A0(\scan_chain.scan_cells[42].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[42].scan_cell.data_in ),
    .S(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_085_));
 sky130_fd_sc_hd__mux2_1 _341_ (.A0(\scan_chain.scan_cells[41].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[40].scan_cell.data_in ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_175_));
 sky130_fd_sc_hd__mux2_1 _342_ (.A0(\scan_chain.scan_cells[41].scan_cell.primary_ff ),
    .A1(_175_),
    .S(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_086_));
 sky130_fd_sc_hd__mux2_1 _343_ (.A0(\scan_chain.scan_cells[41].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[41].scan_cell.data_in ),
    .S(_145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_087_));
 sky130_fd_sc_hd__mux2_1 _344_ (.A0(\scan_chain.scan_cells[40].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[39].scan_cell.data_in ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_176_));
 sky130_fd_sc_hd__mux2_1 _345_ (.A0(\scan_chain.scan_cells[40].scan_cell.primary_ff ),
    .A1(_176_),
    .S(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_088_));
 sky130_fd_sc_hd__mux2_1 _346_ (.A0(\scan_chain.scan_cells[40].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[40].scan_cell.data_in ),
    .S(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_089_));
 sky130_fd_sc_hd__mux2_1 _347_ (.A0(\scan_chain.scan_cells[3].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[2].scan_cell.data_out ),
    .S(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_177_));
 sky130_fd_sc_hd__mux2_1 _348_ (.A0(\scan_chain.scan_cells[3].scan_cell.primary_ff ),
    .A1(_177_),
    .S(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_090_));
 sky130_fd_sc_hd__mux2_1 _349_ (.A0(\scan_chain.scan_cells[39].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[39].scan_cell.data_in ),
    .S(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_091_));
 sky130_fd_sc_hd__mux2_1 _350_ (.A0(\scan_chain.scan_cells[38].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[37].scan_cell.data_in ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_178_));
 sky130_fd_sc_hd__mux2_1 _351_ (.A0(\scan_chain.scan_cells[38].scan_cell.primary_ff ),
    .A1(_178_),
    .S(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_092_));
 sky130_fd_sc_hd__mux2_1 _352_ (.A0(\scan_chain.scan_cells[38].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[38].scan_cell.data_in ),
    .S(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_093_));
 sky130_fd_sc_hd__mux2_1 _353_ (.A0(\scan_chain.scan_cells[37].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[36].scan_cell.data_in ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_179_));
 sky130_fd_sc_hd__mux2_1 _354_ (.A0(\scan_chain.scan_cells[37].scan_cell.primary_ff ),
    .A1(_179_),
    .S(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_094_));
 sky130_fd_sc_hd__mux2_1 _355_ (.A0(\scan_chain.scan_cells[37].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[37].scan_cell.data_in ),
    .S(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_095_));
 sky130_fd_sc_hd__mux2_1 _356_ (.A0(\scan_chain.scan_cells[36].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[35].scan_cell.data_in ),
    .S(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_180_));
 sky130_fd_sc_hd__mux2_1 _357_ (.A0(\scan_chain.scan_cells[36].scan_cell.primary_ff ),
    .A1(_180_),
    .S(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_096_));
 sky130_fd_sc_hd__mux2_1 _358_ (.A0(\scan_chain.scan_cells[36].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[36].scan_cell.data_in ),
    .S(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_097_));
 sky130_fd_sc_hd__mux2_1 _359_ (.A0(\scan_chain.scan_cells[35].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[34].scan_cell.data_in ),
    .S(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_181_));
 sky130_fd_sc_hd__mux2_1 _360_ (.A0(\scan_chain.scan_cells[35].scan_cell.primary_ff ),
    .A1(_181_),
    .S(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_098_));
 sky130_fd_sc_hd__mux2_1 _361_ (.A0(\scan_chain.scan_cells[35].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[35].scan_cell.data_in ),
    .S(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_099_));
 sky130_fd_sc_hd__mux2_1 _362_ (.A0(\scan_chain.scan_cells[34].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[33].scan_cell.data_in ),
    .S(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_182_));
 sky130_fd_sc_hd__mux2_1 _363_ (.A0(\scan_chain.scan_cells[34].scan_cell.primary_ff ),
    .A1(_182_),
    .S(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_100_));
 sky130_fd_sc_hd__mux2_1 _364_ (.A0(\scan_chain.scan_cells[34].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[34].scan_cell.data_in ),
    .S(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_101_));
 sky130_fd_sc_hd__mux2_1 _365_ (.A0(\scan_chain.scan_cells[33].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[32].scan_cell.data_out ),
    .S(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_183_));
 sky130_fd_sc_hd__mux2_1 _366_ (.A0(\scan_chain.scan_cells[33].scan_cell.primary_ff ),
    .A1(_183_),
    .S(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_102_));
 sky130_fd_sc_hd__mux2_1 _367_ (.A0(\scan_chain.scan_cells[33].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[33].scan_cell.data_in ),
    .S(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_103_));
 sky130_fd_sc_hd__mux2_1 _368_ (.A0(\scan_chain.scan_cells[32].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[31].scan_cell.data_out ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_184_));
 sky130_fd_sc_hd__mux2_1 _369_ (.A0(\scan_chain.scan_cells[32].scan_cell.primary_ff ),
    .A1(_184_),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_104_));
 sky130_fd_sc_hd__mux2_1 _370_ (.A0(\dout[32] ),
    .A1(\scan_chain.scan_cells[32].scan_cell.primary_ff ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_185_));
 sky130_fd_sc_hd__mux2_1 _371_ (.A0(\scan_chain.scan_cells[32].scan_cell.data_out ),
    .A1(_185_),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_105_));
 sky130_fd_sc_hd__mux2_1 _372_ (.A0(\scan_chain.scan_cells[31].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[30].scan_cell.data_out ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_186_));
 sky130_fd_sc_hd__mux2_1 _373_ (.A0(\scan_chain.scan_cells[31].scan_cell.primary_ff ),
    .A1(_186_),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_106_));
 sky130_fd_sc_hd__mux2_1 _374_ (.A0(\dout[31] ),
    .A1(\scan_chain.scan_cells[31].scan_cell.primary_ff ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_187_));
 sky130_fd_sc_hd__mux2_1 _375_ (.A0(\scan_chain.scan_cells[31].scan_cell.data_out ),
    .A1(_187_),
    .S(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_107_));
 sky130_fd_sc_hd__mux2_1 _376_ (.A0(\scan_chain.scan_cells[30].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[29].scan_cell.data_out ),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_188_));
 sky130_fd_sc_hd__mux2_1 _377_ (.A0(\scan_chain.scan_cells[30].scan_cell.primary_ff ),
    .A1(_188_),
    .S(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_108_));
 sky130_fd_sc_hd__mux2_1 _378_ (.A0(\dout[30] ),
    .A1(\scan_chain.scan_cells[30].scan_cell.primary_ff ),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_189_));
 sky130_fd_sc_hd__mux2_1 _379_ (.A0(\scan_chain.scan_cells[30].scan_cell.data_out ),
    .A1(_189_),
    .S(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_109_));
 sky130_fd_sc_hd__mux2_1 _380_ (.A0(\scan_chain.scan_cells[2].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[1].scan_cell.data_out ),
    .S(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_190_));
 sky130_fd_sc_hd__mux2_1 _381_ (.A0(\scan_chain.scan_cells[2].scan_cell.primary_ff ),
    .A1(_190_),
    .S(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_110_));
 sky130_fd_sc_hd__mux2_1 _382_ (.A0(\dout[29] ),
    .A1(\scan_chain.scan_cells[29].scan_cell.primary_ff ),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_191_));
 sky130_fd_sc_hd__mux2_1 _383_ (.A0(\scan_chain.scan_cells[29].scan_cell.data_out ),
    .A1(_191_),
    .S(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_111_));
 sky130_fd_sc_hd__mux2_1 _384_ (.A0(\scan_chain.scan_cells[28].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[27].scan_cell.data_out ),
    .S(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_192_));
 sky130_fd_sc_hd__mux2_1 _385_ (.A0(\scan_chain.scan_cells[28].scan_cell.primary_ff ),
    .A1(_192_),
    .S(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_112_));
 sky130_fd_sc_hd__mux2_1 _386_ (.A0(\dout[28] ),
    .A1(\scan_chain.scan_cells[28].scan_cell.primary_ff ),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_193_));
 sky130_fd_sc_hd__mux2_1 _387_ (.A0(\scan_chain.scan_cells[28].scan_cell.data_out ),
    .A1(_193_),
    .S(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_113_));
 sky130_fd_sc_hd__mux2_1 _388_ (.A0(\scan_chain.scan_cells[27].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[26].scan_cell.data_out ),
    .S(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_194_));
 sky130_fd_sc_hd__mux2_1 _389_ (.A0(\scan_chain.scan_cells[27].scan_cell.primary_ff ),
    .A1(_194_),
    .S(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_114_));
 sky130_fd_sc_hd__mux2_1 _390_ (.A0(\dout[27] ),
    .A1(\scan_chain.scan_cells[27].scan_cell.primary_ff ),
    .S(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_195_));
 sky130_fd_sc_hd__mux2_1 _391_ (.A0(\scan_chain.scan_cells[27].scan_cell.data_out ),
    .A1(_195_),
    .S(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_115_));
 sky130_fd_sc_hd__mux2_1 _392_ (.A0(\scan_chain.scan_cells[26].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[25].scan_cell.data_out ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_196_));
 sky130_fd_sc_hd__mux2_1 _393_ (.A0(\scan_chain.scan_cells[26].scan_cell.primary_ff ),
    .A1(_196_),
    .S(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_116_));
 sky130_fd_sc_hd__mux2_1 _394_ (.A0(\dout[26] ),
    .A1(\scan_chain.scan_cells[26].scan_cell.primary_ff ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_197_));
 sky130_fd_sc_hd__mux2_1 _395_ (.A0(\scan_chain.scan_cells[26].scan_cell.data_out ),
    .A1(_197_),
    .S(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_117_));
 sky130_fd_sc_hd__mux2_1 _396_ (.A0(\scan_chain.scan_cells[25].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[24].scan_cell.data_out ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_198_));
 sky130_fd_sc_hd__mux2_1 _397_ (.A0(\scan_chain.scan_cells[25].scan_cell.primary_ff ),
    .A1(_198_),
    .S(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_118_));
 sky130_fd_sc_hd__mux2_1 _398_ (.A0(\dout[25] ),
    .A1(\scan_chain.scan_cells[25].scan_cell.primary_ff ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_199_));
 sky130_fd_sc_hd__mux2_1 _399_ (.A0(\scan_chain.scan_cells[25].scan_cell.data_out ),
    .A1(_199_),
    .S(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_119_));
 sky130_fd_sc_hd__mux2_1 _400_ (.A0(\scan_chain.scan_cells[24].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[23].scan_cell.data_out ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_200_));
 sky130_fd_sc_hd__mux2_1 _401_ (.A0(\scan_chain.scan_cells[24].scan_cell.primary_ff ),
    .A1(_200_),
    .S(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_120_));
 sky130_fd_sc_hd__mux2_1 _402_ (.A0(\dout[24] ),
    .A1(\scan_chain.scan_cells[24].scan_cell.primary_ff ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_201_));
 sky130_fd_sc_hd__mux2_1 _403_ (.A0(\scan_chain.scan_cells[24].scan_cell.data_out ),
    .A1(_201_),
    .S(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_121_));
 sky130_fd_sc_hd__mux2_1 _404_ (.A0(\scan_chain.scan_cells[23].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[22].scan_cell.data_out ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_202_));
 sky130_fd_sc_hd__mux2_1 _405_ (.A0(\scan_chain.scan_cells[23].scan_cell.primary_ff ),
    .A1(_202_),
    .S(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_122_));
 sky130_fd_sc_hd__mux2_1 _406_ (.A0(\dout[23] ),
    .A1(\scan_chain.scan_cells[23].scan_cell.primary_ff ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_203_));
 sky130_fd_sc_hd__mux2_1 _407_ (.A0(\scan_chain.scan_cells[23].scan_cell.data_out ),
    .A1(_203_),
    .S(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_123_));
 sky130_fd_sc_hd__mux2_1 _408_ (.A0(\scan_chain.scan_cells[22].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[21].scan_cell.data_out ),
    .S(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_204_));
 sky130_fd_sc_hd__mux2_1 _409_ (.A0(\scan_chain.scan_cells[22].scan_cell.primary_ff ),
    .A1(_204_),
    .S(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_124_));
 sky130_fd_sc_hd__mux2_1 _410_ (.A0(\dout[22] ),
    .A1(\scan_chain.scan_cells[22].scan_cell.primary_ff ),
    .S(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_205_));
 sky130_fd_sc_hd__mux2_1 _411_ (.A0(\scan_chain.scan_cells[22].scan_cell.data_out ),
    .A1(_205_),
    .S(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_125_));
 sky130_fd_sc_hd__mux2_1 _412_ (.A0(\scan_chain.scan_cells[21].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[20].scan_cell.data_out ),
    .S(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_206_));
 sky130_fd_sc_hd__mux2_1 _413_ (.A0(\scan_chain.scan_cells[21].scan_cell.primary_ff ),
    .A1(_206_),
    .S(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_126_));
 sky130_fd_sc_hd__mux2_1 _414_ (.A0(\dout[21] ),
    .A1(\scan_chain.scan_cells[21].scan_cell.primary_ff ),
    .S(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_207_));
 sky130_fd_sc_hd__mux2_1 _415_ (.A0(\scan_chain.scan_cells[21].scan_cell.data_out ),
    .A1(_207_),
    .S(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_127_));
 sky130_fd_sc_hd__mux2_1 _416_ (.A0(\scan_chain.scan_cells[20].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[19].scan_cell.data_out ),
    .S(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_208_));
 sky130_fd_sc_hd__mux2_1 _417_ (.A0(\scan_chain.scan_cells[20].scan_cell.primary_ff ),
    .A1(_208_),
    .S(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_128_));
 sky130_fd_sc_hd__mux2_1 _418_ (.A0(\dout[20] ),
    .A1(\scan_chain.scan_cells[20].scan_cell.primary_ff ),
    .S(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_209_));
 sky130_fd_sc_hd__mux2_1 _419_ (.A0(\scan_chain.scan_cells[20].scan_cell.data_out ),
    .A1(_209_),
    .S(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_129_));
 sky130_fd_sc_hd__mux2_1 _420_ (.A0(\scan_chain.scan_cells[1].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[0].scan_cell.data_out ),
    .S(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_210_));
 sky130_fd_sc_hd__mux2_1 _421_ (.A0(\scan_chain.scan_cells[1].scan_cell.primary_ff ),
    .A1(_210_),
    .S(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_130_));
 sky130_fd_sc_hd__mux2_1 _422_ (.A0(\dout[19] ),
    .A1(\scan_chain.scan_cells[19].scan_cell.primary_ff ),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_211_));
 sky130_fd_sc_hd__mux2_1 _423_ (.A0(\scan_chain.scan_cells[19].scan_cell.data_out ),
    .A1(_211_),
    .S(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_131_));
 sky130_fd_sc_hd__mux2_1 _424_ (.A0(\scan_chain.scan_cells[18].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[17].scan_cell.data_out ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_212_));
 sky130_fd_sc_hd__mux2_1 _425_ (.A0(\scan_chain.scan_cells[18].scan_cell.primary_ff ),
    .A1(_212_),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_132_));
 sky130_fd_sc_hd__mux2_1 _426_ (.A0(\dout[18] ),
    .A1(\scan_chain.scan_cells[18].scan_cell.primary_ff ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_213_));
 sky130_fd_sc_hd__mux2_1 _427_ (.A0(\scan_chain.scan_cells[18].scan_cell.data_out ),
    .A1(_213_),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_133_));
 sky130_fd_sc_hd__mux2_1 _428_ (.A0(\scan_chain.scan_cells[17].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[16].scan_cell.data_out ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_214_));
 sky130_fd_sc_hd__mux2_1 _429_ (.A0(\scan_chain.scan_cells[17].scan_cell.primary_ff ),
    .A1(_214_),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_134_));
 sky130_fd_sc_hd__mux2_1 _430_ (.A0(\dout[17] ),
    .A1(\scan_chain.scan_cells[17].scan_cell.primary_ff ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_215_));
 sky130_fd_sc_hd__mux2_1 _431_ (.A0(\scan_chain.scan_cells[17].scan_cell.data_out ),
    .A1(_215_),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_135_));
 sky130_fd_sc_hd__mux2_1 _432_ (.A0(\scan_chain.scan_cells[16].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[15].scan_cell.data_out ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_216_));
 sky130_fd_sc_hd__mux2_1 _433_ (.A0(\scan_chain.scan_cells[16].scan_cell.primary_ff ),
    .A1(_216_),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_136_));
 sky130_fd_sc_hd__mux2_1 _434_ (.A0(\dout[16] ),
    .A1(\scan_chain.scan_cells[16].scan_cell.primary_ff ),
    .S(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_217_));
 sky130_fd_sc_hd__mux2_1 _435_ (.A0(\scan_chain.scan_cells[16].scan_cell.data_out ),
    .A1(_217_),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_137_));
 sky130_fd_sc_hd__mux2_1 _436_ (.A0(\scan_chain.scan_cells[15].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[14].scan_cell.data_out ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_218_));
 sky130_fd_sc_hd__mux2_1 _437_ (.A0(\scan_chain.scan_cells[15].scan_cell.primary_ff ),
    .A1(_218_),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_138_));
 sky130_fd_sc_hd__mux2_1 _438_ (.A0(\dout[15] ),
    .A1(\scan_chain.scan_cells[15].scan_cell.primary_ff ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_219_));
 sky130_fd_sc_hd__mux2_1 _439_ (.A0(\scan_chain.scan_cells[15].scan_cell.data_out ),
    .A1(_219_),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_139_));
 sky130_fd_sc_hd__mux2_1 _440_ (.A0(\scan_chain.scan_cells[14].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[13].scan_cell.data_out ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_220_));
 sky130_fd_sc_hd__mux2_1 _441_ (.A0(\scan_chain.scan_cells[14].scan_cell.primary_ff ),
    .A1(_220_),
    .S(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_140_));
 sky130_fd_sc_hd__mux2_1 _442_ (.A0(\dout[14] ),
    .A1(\scan_chain.scan_cells[14].scan_cell.primary_ff ),
    .S(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_221_));
 sky130_fd_sc_hd__mux2_1 _443_ (.A0(\scan_chain.scan_cells[14].scan_cell.data_out ),
    .A1(_221_),
    .S(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_141_));
 sky130_fd_sc_hd__mux2_1 _444_ (.A0(\scan_chain.scan_cells[13].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[12].scan_cell.data_out ),
    .S(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_222_));
 sky130_fd_sc_hd__mux2_1 _445_ (.A0(\scan_chain.scan_cells[13].scan_cell.primary_ff ),
    .A1(_222_),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_142_));
 sky130_fd_sc_hd__mux2_1 _446_ (.A0(\dout[13] ),
    .A1(\scan_chain.scan_cells[13].scan_cell.primary_ff ),
    .S(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_223_));
 sky130_fd_sc_hd__mux2_1 _447_ (.A0(\scan_chain.scan_cells[13].scan_cell.data_out ),
    .A1(_223_),
    .S(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_143_));
 sky130_fd_sc_hd__mux2_1 _448_ (.A0(\scan_chain.scan_cells[12].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[11].scan_cell.data_out ),
    .S(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_224_));
 sky130_fd_sc_hd__mux2_1 _449_ (.A0(\scan_chain.scan_cells[12].scan_cell.primary_ff ),
    .A1(_224_),
    .S(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_000_));
 sky130_fd_sc_hd__mux2_1 _450_ (.A0(\dout[12] ),
    .A1(\scan_chain.scan_cells[12].scan_cell.primary_ff ),
    .S(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_225_));
 sky130_fd_sc_hd__mux2_1 _451_ (.A0(\scan_chain.scan_cells[12].scan_cell.data_out ),
    .A1(_225_),
    .S(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _452_ (.A0(\scan_chain.scan_cells[11].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[10].scan_cell.data_out ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_226_));
 sky130_fd_sc_hd__mux2_1 _453_ (.A0(\scan_chain.scan_cells[11].scan_cell.primary_ff ),
    .A1(_226_),
    .S(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _454_ (.A0(\dout[11] ),
    .A1(\scan_chain.scan_cells[11].scan_cell.primary_ff ),
    .S(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_227_));
 sky130_fd_sc_hd__mux2_1 _455_ (.A0(\scan_chain.scan_cells[11].scan_cell.data_out ),
    .A1(_227_),
    .S(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _456_ (.A0(\scan_chain.scan_cells[10].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[10].scan_cell.scan_in ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_228_));
 sky130_fd_sc_hd__mux2_1 _457_ (.A0(\scan_chain.scan_cells[10].scan_cell.primary_ff ),
    .A1(_228_),
    .S(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _458_ (.A0(\dout[10] ),
    .A1(\scan_chain.scan_cells[10].scan_cell.primary_ff ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_229_));
 sky130_fd_sc_hd__mux2_1 _459_ (.A0(\scan_chain.scan_cells[10].scan_cell.data_out ),
    .A1(_229_),
    .S(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _460_ (.A0(\scan_chain.scan_cells[0].scan_cell.data_out ),
    .A1(net2),
    .S(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_230_));
 sky130_fd_sc_hd__mux2_1 _461_ (.A0(\scan_chain.scan_cells[0].scan_cell.primary_ff ),
    .A1(_230_),
    .S(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _462_ (.A0(\dout[9] ),
    .A1(\scan_chain.scan_cells[9].scan_cell.primary_ff ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_231_));
 sky130_fd_sc_hd__mux2_1 _463_ (.A0(\scan_chain.scan_cells[10].scan_cell.scan_in ),
    .A1(_231_),
    .S(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _464_ (.A0(\scan_chain.scan_cells[8].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[7].scan_cell.data_out ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_232_));
 sky130_fd_sc_hd__mux2_1 _465_ (.A0(\scan_chain.scan_cells[8].scan_cell.primary_ff ),
    .A1(_232_),
    .S(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _466_ (.A0(\dout[8] ),
    .A1(\scan_chain.scan_cells[8].scan_cell.primary_ff ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_233_));
 sky130_fd_sc_hd__mux2_1 _467_ (.A0(\scan_chain.scan_cells[8].scan_cell.data_out ),
    .A1(_233_),
    .S(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _468_ (.A0(\scan_chain.scan_cells[7].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[6].scan_cell.data_out ),
    .S(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_234_));
 sky130_fd_sc_hd__mux2_1 _469_ (.A0(\scan_chain.scan_cells[7].scan_cell.primary_ff ),
    .A1(_234_),
    .S(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _470_ (.A0(\dout[7] ),
    .A1(\scan_chain.scan_cells[7].scan_cell.primary_ff ),
    .S(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_235_));
 sky130_fd_sc_hd__mux2_1 _471_ (.A0(\scan_chain.scan_cells[7].scan_cell.data_out ),
    .A1(_235_),
    .S(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _472_ (.A0(\scan_chain.scan_cells[71].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[70].scan_cell.data_in ),
    .S(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_236_));
 sky130_fd_sc_hd__mux2_1 _473_ (.A0(\scan_chain.scan_cells[71].scan_cell.primary_ff ),
    .A1(_236_),
    .S(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _474_ (.A0(\dout[6] ),
    .A1(\scan_chain.scan_cells[6].scan_cell.primary_ff ),
    .S(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_237_));
 sky130_fd_sc_hd__mux2_1 _475_ (.A0(\scan_chain.scan_cells[6].scan_cell.data_out ),
    .A1(_237_),
    .S(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _476_ (.A0(\scan_chain.scan_cells[69].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[68].scan_cell.data_in ),
    .S(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_238_));
 sky130_fd_sc_hd__mux2_1 _477_ (.A0(\scan_chain.scan_cells[69].scan_cell.primary_ff ),
    .A1(_238_),
    .S(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _478_ (.A0(\dout[5] ),
    .A1(\scan_chain.scan_cells[5].scan_cell.primary_ff ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_239_));
 sky130_fd_sc_hd__mux2_1 _479_ (.A0(\scan_chain.scan_cells[5].scan_cell.data_out ),
    .A1(_239_),
    .S(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _480_ (.A0(\scan_chain.scan_cells[59].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[58].scan_cell.data_in ),
    .S(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_240_));
 sky130_fd_sc_hd__mux2_1 _481_ (.A0(\scan_chain.scan_cells[59].scan_cell.primary_ff ),
    .A1(_240_),
    .S(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _482_ (.A0(\dout[4] ),
    .A1(\scan_chain.scan_cells[4].scan_cell.primary_ff ),
    .S(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_241_));
 sky130_fd_sc_hd__mux2_1 _483_ (.A0(\scan_chain.scan_cells[4].scan_cell.data_out ),
    .A1(_241_),
    .S(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _484_ (.A0(\scan_chain.scan_cells[49].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[48].scan_cell.data_in ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_242_));
 sky130_fd_sc_hd__mux2_1 _485_ (.A0(\scan_chain.scan_cells[49].scan_cell.primary_ff ),
    .A1(_242_),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_018_));
 sky130_fd_sc_hd__mux2_1 _486_ (.A0(\dout[3] ),
    .A1(\scan_chain.scan_cells[3].scan_cell.primary_ff ),
    .S(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_243_));
 sky130_fd_sc_hd__mux2_1 _487_ (.A0(\scan_chain.scan_cells[3].scan_cell.data_out ),
    .A1(_243_),
    .S(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_019_));
 sky130_fd_sc_hd__mux2_1 _488_ (.A0(\scan_chain.scan_cells[39].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[38].scan_cell.data_in ),
    .S(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_244_));
 sky130_fd_sc_hd__mux2_1 _489_ (.A0(\scan_chain.scan_cells[39].scan_cell.primary_ff ),
    .A1(_244_),
    .S(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_020_));
 sky130_fd_sc_hd__mux2_1 _490_ (.A0(\dout[2] ),
    .A1(\scan_chain.scan_cells[2].scan_cell.primary_ff ),
    .S(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_245_));
 sky130_fd_sc_hd__mux2_1 _491_ (.A0(\scan_chain.scan_cells[2].scan_cell.data_out ),
    .A1(_245_),
    .S(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _492_ (.A0(\scan_chain.scan_cells[29].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[28].scan_cell.data_out ),
    .S(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_246_));
 sky130_fd_sc_hd__mux2_1 _493_ (.A0(\scan_chain.scan_cells[29].scan_cell.primary_ff ),
    .A1(_246_),
    .S(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_022_));
 sky130_fd_sc_hd__mux2_1 _494_ (.A0(\dout[1] ),
    .A1(\scan_chain.scan_cells[1].scan_cell.primary_ff ),
    .S(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_247_));
 sky130_fd_sc_hd__mux2_1 _495_ (.A0(\scan_chain.scan_cells[1].scan_cell.data_out ),
    .A1(_247_),
    .S(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_023_));
 sky130_fd_sc_hd__mux2_1 _496_ (.A0(\scan_chain.scan_cells[19].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[18].scan_cell.data_out ),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_248_));
 sky130_fd_sc_hd__mux2_1 _497_ (.A0(\scan_chain.scan_cells[19].scan_cell.primary_ff ),
    .A1(_248_),
    .S(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _498_ (.A0(\dout[0] ),
    .A1(\scan_chain.scan_cells[0].scan_cell.primary_ff ),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_249_));
 sky130_fd_sc_hd__mux2_1 _499_ (.A0(\scan_chain.scan_cells[0].scan_cell.data_out ),
    .A1(_249_),
    .S(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_025_));
 sky130_fd_sc_hd__dfrtp_1 _500_ (.CLK(clknet_3_0__leaf_ui_in[3]),
    .D(_026_),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[9].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _501_ (.CLK(clknet_3_2__leaf_ui_in[4]),
    .D(_027_),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[71].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _502_ (.CLK(clknet_3_2__leaf_ui_in[3]),
    .D(_028_),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[70].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _503_ (.CLK(clknet_3_2__leaf_ui_in[4]),
    .D(_029_),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[70].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _504_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_030_),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[6].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _505_ (.CLK(clknet_3_2__leaf_ui_in[4]),
    .D(_031_),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[69].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _506_ (.CLK(clknet_3_2__leaf_ui_in[3]),
    .D(_032_),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[68].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _507_ (.CLK(clknet_3_2__leaf_ui_in[4]),
    .D(_033_),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[68].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _508_ (.CLK(clknet_3_2__leaf_ui_in[3]),
    .D(_034_),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[67].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _509_ (.CLK(clknet_3_2__leaf_ui_in[4]),
    .D(_035_),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[67].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _510_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_036_),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[66].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _511_ (.CLK(clknet_3_2__leaf_ui_in[4]),
    .D(_037_),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[66].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _512_ (.CLK(clknet_3_7__leaf_ui_in[3]),
    .D(_038_),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[65].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _513_ (.CLK(clknet_3_4__leaf_ui_in[4]),
    .D(_039_),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[65].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _514_ (.CLK(clknet_3_7__leaf_ui_in[3]),
    .D(_040_),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[64].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _515_ (.CLK(clknet_3_4__leaf_ui_in[4]),
    .D(_041_),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[64].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _516_ (.CLK(clknet_3_4__leaf_ui_in[3]),
    .D(_042_),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[63].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _517_ (.CLK(clknet_3_4__leaf_ui_in[4]),
    .D(_043_),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[63].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _518_ (.CLK(clknet_3_4__leaf_ui_in[3]),
    .D(_044_),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[62].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _519_ (.CLK(clknet_3_4__leaf_ui_in[4]),
    .D(_045_),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[62].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _520_ (.CLK(clknet_3_7__leaf_ui_in[3]),
    .D(_046_),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[61].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _521_ (.CLK(clknet_3_7__leaf_ui_in[4]),
    .D(_047_),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[61].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _522_ (.CLK(clknet_3_7__leaf_ui_in[3]),
    .D(_048_),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[60].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _523_ (.CLK(clknet_3_7__leaf_ui_in[4]),
    .D(_049_),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[60].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _524_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_050_),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[5].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _525_ (.CLK(clknet_3_7__leaf_ui_in[4]),
    .D(_051_),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[59].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _526_ (.CLK(clknet_3_4__leaf_ui_in[3]),
    .D(_052_),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[58].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _527_ (.CLK(clknet_3_7__leaf_ui_in[4]),
    .D(_053_),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[58].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _528_ (.CLK(clknet_3_7__leaf_ui_in[3]),
    .D(_054_),
    .RESET_B(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[57].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_2 _529_ (.CLK(clknet_3_7__leaf_ui_in[4]),
    .D(_055_),
    .RESET_B(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[57].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _530_ (.CLK(clknet_3_7__leaf_ui_in[3]),
    .D(_056_),
    .RESET_B(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[56].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _531_ (.CLK(clknet_3_7__leaf_ui_in[4]),
    .D(_057_),
    .RESET_B(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[56].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _532_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_058_),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[55].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_2 _533_ (.CLK(clknet_3_7__leaf_ui_in[4]),
    .D(_059_),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[55].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _534_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_060_),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[54].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_2 _535_ (.CLK(clknet_3_7__leaf_ui_in[4]),
    .D(_061_),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[54].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _536_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_062_),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[53].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_2 _537_ (.CLK(clknet_3_7__leaf_ui_in[4]),
    .D(_063_),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[53].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _538_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_064_),
    .RESET_B(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[52].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_2 _539_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_065_),
    .RESET_B(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[52].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _540_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_066_),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[51].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_2 _541_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_067_),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[51].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _542_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_068_),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[50].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _543_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_069_),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[50].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _544_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_070_),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[4].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _545_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_071_),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[49].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _546_ (.CLK(clknet_3_1__leaf_ui_in[3]),
    .D(_072_),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[48].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _547_ (.CLK(clknet_3_1__leaf_ui_in[4]),
    .D(_073_),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[48].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _548_ (.CLK(clknet_3_1__leaf_ui_in[3]),
    .D(_074_),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[47].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _549_ (.CLK(clknet_3_1__leaf_ui_in[4]),
    .D(_075_),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[47].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _550_ (.CLK(clknet_3_0__leaf_ui_in[3]),
    .D(_076_),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[46].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _551_ (.CLK(clknet_3_0__leaf_ui_in[4]),
    .D(_077_),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[46].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _552_ (.CLK(clknet_3_0__leaf_ui_in[3]),
    .D(_078_),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[45].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _553_ (.CLK(clknet_3_0__leaf_ui_in[4]),
    .D(_079_),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[45].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _554_ (.CLK(clknet_3_0__leaf_ui_in[3]),
    .D(_080_),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[44].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _555_ (.CLK(clknet_3_0__leaf_ui_in[4]),
    .D(_081_),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[44].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _556_ (.CLK(clknet_3_0__leaf_ui_in[3]),
    .D(_082_),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[43].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _557_ (.CLK(clknet_3_0__leaf_ui_in[4]),
    .D(_083_),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[43].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _558_ (.CLK(clknet_3_2__leaf_ui_in[3]),
    .D(_084_),
    .RESET_B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[42].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _559_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_085_),
    .RESET_B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[42].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _560_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_086_),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[41].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _561_ (.CLK(clknet_3_0__leaf_ui_in[4]),
    .D(_087_),
    .RESET_B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[41].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _562_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_088_),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[40].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _563_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_089_),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[40].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _564_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_090_),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[3].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _565_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_091_),
    .RESET_B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[39].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _566_ (.CLK(clknet_3_2__leaf_ui_in[3]),
    .D(_092_),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[38].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _567_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_093_),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[38].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _568_ (.CLK(clknet_3_2__leaf_ui_in[3]),
    .D(_094_),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[37].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _569_ (.CLK(clknet_3_2__leaf_ui_in[4]),
    .D(_095_),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[37].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _570_ (.CLK(clknet_3_2__leaf_ui_in[3]),
    .D(_096_),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[36].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _571_ (.CLK(clknet_3_2__leaf_ui_in[4]),
    .D(_097_),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[36].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _572_ (.CLK(clknet_3_2__leaf_ui_in[3]),
    .D(_098_),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[35].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_2 _573_ (.CLK(clknet_3_2__leaf_ui_in[4]),
    .D(_099_),
    .RESET_B(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[35].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _574_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_100_),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[34].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_2 _575_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_101_),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[34].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _576_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_102_),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[33].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_2 _577_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_103_),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[33].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _578_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_104_),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[32].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _579_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_105_),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[32].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _580_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_106_),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[31].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _581_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_107_),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[31].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _582_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_108_),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[30].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _583_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_109_),
    .RESET_B(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[30].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _584_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_110_),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[2].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _585_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_111_),
    .RESET_B(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[29].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _586_ (.CLK(clknet_3_4__leaf_ui_in[3]),
    .D(_112_),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[28].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _587_ (.CLK(clknet_3_7__leaf_ui_in[4]),
    .D(_113_),
    .RESET_B(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[28].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _588_ (.CLK(clknet_3_4__leaf_ui_in[3]),
    .D(_114_),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[27].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _589_ (.CLK(clknet_3_4__leaf_ui_in[4]),
    .D(_115_),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[27].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _590_ (.CLK(clknet_3_5__leaf_ui_in[3]),
    .D(_116_),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[26].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _591_ (.CLK(clknet_3_5__leaf_ui_in[4]),
    .D(_117_),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[26].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _592_ (.CLK(clknet_3_5__leaf_ui_in[3]),
    .D(_118_),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[25].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _593_ (.CLK(clknet_3_5__leaf_ui_in[4]),
    .D(_119_),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[25].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _594_ (.CLK(clknet_3_5__leaf_ui_in[3]),
    .D(_120_),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[24].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _595_ (.CLK(clknet_3_5__leaf_ui_in[4]),
    .D(_121_),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[24].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _596_ (.CLK(clknet_3_5__leaf_ui_in[3]),
    .D(_122_),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[23].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _597_ (.CLK(clknet_3_5__leaf_ui_in[4]),
    .D(_123_),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[23].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _598_ (.CLK(clknet_3_5__leaf_ui_in[3]),
    .D(_124_),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[22].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _599_ (.CLK(clknet_3_5__leaf_ui_in[4]),
    .D(_125_),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[22].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _600_ (.CLK(clknet_3_4__leaf_ui_in[3]),
    .D(_126_),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[21].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _601_ (.CLK(clknet_3_4__leaf_ui_in[4]),
    .D(_127_),
    .RESET_B(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[21].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _602_ (.CLK(clknet_3_7__leaf_ui_in[3]),
    .D(_128_),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[20].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _603_ (.CLK(clknet_3_4__leaf_ui_in[4]),
    .D(_129_),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[20].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _604_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_130_),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[1].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _605_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_131_),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[19].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _606_ (.CLK(clknet_3_1__leaf_ui_in[3]),
    .D(_132_),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[18].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _607_ (.CLK(clknet_3_1__leaf_ui_in[4]),
    .D(_133_),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[18].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _608_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_134_),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[17].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _609_ (.CLK(clknet_3_1__leaf_ui_in[4]),
    .D(_135_),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[17].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _610_ (.CLK(clknet_3_1__leaf_ui_in[3]),
    .D(_136_),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[16].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _611_ (.CLK(clknet_3_1__leaf_ui_in[4]),
    .D(_137_),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[16].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _612_ (.CLK(clknet_3_1__leaf_ui_in[3]),
    .D(_138_),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[15].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _613_ (.CLK(clknet_3_1__leaf_ui_in[4]),
    .D(_139_),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[15].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _614_ (.CLK(clknet_3_1__leaf_ui_in[3]),
    .D(_140_),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[14].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _615_ (.CLK(clknet_3_0__leaf_ui_in[4]),
    .D(_141_),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[14].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _616_ (.CLK(clknet_3_1__leaf_ui_in[3]),
    .D(_142_),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[13].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _617_ (.CLK(clknet_3_1__leaf_ui_in[4]),
    .D(_143_),
    .RESET_B(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[13].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _618_ (.CLK(clknet_3_5__leaf_ui_in[3]),
    .D(_000_),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[12].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _619_ (.CLK(clknet_3_5__leaf_ui_in[4]),
    .D(_001_),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[12].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _620_ (.CLK(clknet_3_5__leaf_ui_in[3]),
    .D(_002_),
    .RESET_B(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[11].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _621_ (.CLK(clknet_3_5__leaf_ui_in[4]),
    .D(_003_),
    .RESET_B(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[11].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _622_ (.CLK(clknet_3_0__leaf_ui_in[3]),
    .D(_004_),
    .RESET_B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[10].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _623_ (.CLK(clknet_3_0__leaf_ui_in[4]),
    .D(_005_),
    .RESET_B(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[10].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _624_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_006_),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[0].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _625_ (.CLK(clknet_3_0__leaf_ui_in[4]),
    .D(_007_),
    .RESET_B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[10].scan_cell.scan_in ));
 sky130_fd_sc_hd__dfrtp_1 _626_ (.CLK(clknet_3_0__leaf_ui_in[3]),
    .D(_008_),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[8].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _627_ (.CLK(clknet_3_0__leaf_ui_in[4]),
    .D(_009_),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[8].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _628_ (.CLK(clknet_3_0__leaf_ui_in[3]),
    .D(_010_),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[7].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _629_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_011_),
    .RESET_B(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[7].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _630_ (.CLK(clknet_3_2__leaf_ui_in[3]),
    .D(_012_),
    .RESET_B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[71].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _631_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_013_),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[6].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _632_ (.CLK(clknet_3_2__leaf_ui_in[3]),
    .D(_014_),
    .RESET_B(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[69].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _633_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_015_),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[5].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _634_ (.CLK(clknet_3_7__leaf_ui_in[3]),
    .D(_016_),
    .RESET_B(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[59].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _635_ (.CLK(clknet_3_2__leaf_ui_in[4]),
    .D(_017_),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[4].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _636_ (.CLK(clknet_3_1__leaf_ui_in[3]),
    .D(_018_),
    .RESET_B(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[49].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _637_ (.CLK(clknet_3_2__leaf_ui_in[4]),
    .D(_019_),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[3].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _638_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_020_),
    .RESET_B(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[39].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _639_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_021_),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[2].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _640_ (.CLK(clknet_3_7__leaf_ui_in[3]),
    .D(_022_),
    .RESET_B(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[29].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _641_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_023_),
    .RESET_B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[1].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _642_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_024_),
    .RESET_B(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[19].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _643_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_025_),
    .RESET_B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\scan_chain.scan_cells[0].scan_cell.data_out ));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net57));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net58));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net59));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net60));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net61));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net62));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net63));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net64));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net65));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net66));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net67));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net68));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net69));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net70));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net71));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net72));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net73));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net74));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net75));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net76));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net77));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_ui_in[3]  (.A(ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_ui_in[3]));
 sky130_fd_sc_hd__buf_2 _666_ (.A(\scan_chain.scan_cells[71].scan_cell.data_in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__buf_2 _667_ (.A(\scan_chain.scan_cells[0].scan_cell.data_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[1]));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_2_Left_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_2_Left_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_2_Left_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_2_Left_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_2_Left_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_2_Left_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_2_Left_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_2_Left_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_2_Left_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Left_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Left_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Left_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Left_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Left_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Left_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Left_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Left_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Left_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Left_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Left_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Left_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Left_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Left_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Left_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Left_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Left_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Left_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Left_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Left_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Left_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Left_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Left_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Left_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Left_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Left_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Left_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Left_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Left_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Left_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Left_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Left_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Left_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Left_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Left_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Left_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Left_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Left_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Left_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Left_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Left_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Left_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Left_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Left_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Left_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Left_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Left_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Left_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Left_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Left_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Left_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Left_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Left_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Left_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Left_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Left_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Left_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_2_Left_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_2_Right_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_2_Right_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_2_Right_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_2_Right_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_2_Right_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_2_Right_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_2_Right_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_2_Right_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_2_Right_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Right_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Right_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Right_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Right_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Right_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Right_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Right_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Right_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Right_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Right_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Right_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Right_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Right_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Right_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Right_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Right_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Right_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Right_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Right_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Right_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Right_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Right_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Right_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Right_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Right_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Right_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Right_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Right_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Right_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Right_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Right_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Right_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Right_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Right_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Right_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Right_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Right_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Right_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Right_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Right_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Right_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Right_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Right_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Right_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Right_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Right_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Right_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Right_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Right_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Right_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Right_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Right_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Right_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Right_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Right_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Right_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Right_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_2_Right_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(ui_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 fanout5 (.A(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 fanout6 (.A(_145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 fanout7 (.A(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 fanout8 (.A(_145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 fanout9 (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 fanout10 (.A(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 fanout11 (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 fanout12 (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 fanout13 (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 fanout14 (.A(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 fanout15 (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 fanout16 (.A(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__buf_4 fanout17 (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 fanout18 (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 fanout19 (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__buf_2 fanout20 (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 fanout21 (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__buf_2 fanout22 (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__buf_4 fanout23 (.A(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 fanout24 (.A(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__buf_2 fanout25 (.A(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 fanout26 (.A(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 fanout27 (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 fanout28 (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
 sky130_fd_sc_hd__buf_2 fanout29 (.A(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 fanout30 (.A(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 fanout31 (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net31));
 sky130_fd_sc_hd__buf_2 fanout32 (.A(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 fanout33 (.A(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 fanout34 (.A(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net34));
 sky130_fd_sc_hd__buf_2 fanout35 (.A(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net35));
 sky130_fd_sc_hd__buf_4 fanout36 (.A(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 fanout37 (.A(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 fanout38 (.A(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net38));
 sky130_fd_sc_hd__buf_2 fanout39 (.A(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_4 fanout40 (.A(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net40));
 sky130_fd_sc_hd__buf_2 fanout41 (.A(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net42));
 sky130_fd_sc_hd__buf_2 fanout43 (.A(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 fanout44 (.A(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net44));
 sky130_fd_sc_hd__buf_2 fanout45 (.A(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 fanout46 (.A(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 fanout47 (.A(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__buf_2 fanout48 (.A(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 fanout49 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 fanout50 (.A(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 fanout51 (.A(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 fanout52 (.A(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net52));
 sky130_fd_sc_hd__buf_2 fanout53 (.A(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net53));
 sky130_fd_sc_hd__buf_4 fanout54 (.A(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 fanout55 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net55));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net56));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_0__f_ui_in[3]  (.A(clknet_0_ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_0__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_1__f_ui_in[3]  (.A(clknet_0_ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_1__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_2__f_ui_in[3]  (.A(clknet_0_ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_2__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_3__f_ui_in[3]  (.A(clknet_0_ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_3__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_4__f_ui_in[3]  (.A(clknet_0_ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_4__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_5__f_ui_in[3]  (.A(clknet_0_ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_5__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_6__f_ui_in[3]  (.A(clknet_0_ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_6__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_7__f_ui_in[3]  (.A(clknet_0_ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_7__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkinvlp_4 clkload0 (.A(clknet_3_0__leaf_ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinvlp_4 clkload1 (.A(clknet_3_1__leaf_ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_2 clkload2 (.A(clknet_3_2__leaf_ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_6 clkload3 (.A(clknet_3_4__leaf_ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_4 clkload4 (.A(clknet_3_5__leaf_ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_8 clkload5 (.A(clknet_3_6__leaf_ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__bufinv_16 clkload6 (.A(clknet_3_7__leaf_ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_ui_in[4]  (.A(ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_ui_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_0__f_ui_in[4]  (.A(clknet_0_ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_0__leaf_ui_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_1__f_ui_in[4]  (.A(clknet_0_ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_1__leaf_ui_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_2__f_ui_in[4]  (.A(clknet_0_ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_2__leaf_ui_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_3__f_ui_in[4]  (.A(clknet_0_ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_3__leaf_ui_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_4__f_ui_in[4]  (.A(clknet_0_ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_4__leaf_ui_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_5__f_ui_in[4]  (.A(clknet_0_ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_5__leaf_ui_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_6__f_ui_in[4]  (.A(clknet_0_ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_6__leaf_ui_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_7__f_ui_in[4]  (.A(clknet_0_ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_7__leaf_ui_in[4]));
 sky130_fd_sc_hd__clkinv_2 clkload7 (.A(clknet_3_0__leaf_ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinvlp_4 clkload8 (.A(clknet_3_1__leaf_ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload9 (.A(clknet_3_2__leaf_ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinvlp_4 clkload10 (.A(clknet_3_4__leaf_ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinvlp_4 clkload11 (.A(clknet_3_5__leaf_ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_2 clkload12 (.A(clknet_3_6__leaf_ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_8 clkload13 (.A(clknet_3_7__leaf_ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 assign uio_oe[0] = net56;
 assign uio_oe[1] = net57;
 assign uio_oe[2] = net58;
 assign uio_oe[3] = net59;
 assign uio_oe[4] = net60;
 assign uio_oe[5] = net61;
 assign uio_oe[6] = net62;
 assign uio_oe[7] = net63;
 assign uio_out[0] = net64;
 assign uio_out[1] = net65;
 assign uio_out[2] = net66;
 assign uio_out[3] = net67;
 assign uio_out[4] = net68;
 assign uio_out[5] = net69;
 assign uio_out[6] = net70;
 assign uio_out[7] = net71;
 assign uo_out[2] = net72;
 assign uo_out[3] = net73;
 assign uo_out[4] = net74;
 assign uo_out[5] = net75;
 assign uo_out[6] = net76;
 assign uo_out[7] = net77;
endmodule
