VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_sram_256B_1rw_32x64
  CLASS BLOCK ;
  FOREIGN sky130_sram_256B_1rw_32x64 ;
  ORIGIN 0.000 0.000 ;
  SIZE 310.680 BY 167.570 ;
  SYMMETRY X Y R90 ;
  PIN din0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 100.540 0.000 100.920 0.380 ;
    END
  END din0[0]
  PIN din0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 106.380 0.000 106.760 0.380 ;
    END
  END din0[1]
  PIN din0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 112.220 0.000 112.600 0.380 ;
    END
  END din0[2]
  PIN din0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 118.060 0.000 118.440 0.380 ;
    END
  END din0[3]
  PIN din0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 123.900 0.000 124.280 0.380 ;
    END
  END din0[4]
  PIN din0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 129.740 0.000 130.120 0.380 ;
    END
  END din0[5]
  PIN din0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 135.580 0.000 135.960 0.380 ;
    END
  END din0[6]
  PIN din0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 141.420 0.000 141.800 0.380 ;
    END
  END din0[7]
  PIN din0[8]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 147.260 0.000 147.640 0.380 ;
    END
  END din0[8]
  PIN din0[9]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 153.100 0.000 153.480 0.380 ;
    END
  END din0[9]
  PIN din0[10]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 158.940 0.000 159.320 0.380 ;
    END
  END din0[10]
  PIN din0[11]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 164.780 0.000 165.160 0.380 ;
    END
  END din0[11]
  PIN din0[12]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 170.620 0.000 171.000 0.380 ;
    END
  END din0[12]
  PIN din0[13]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 176.460 0.000 176.840 0.380 ;
    END
  END din0[13]
  PIN din0[14]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 182.300 0.000 182.680 0.380 ;
    END
  END din0[14]
  PIN din0[15]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 188.140 0.000 188.520 0.380 ;
    END
  END din0[15]
  PIN din0[16]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 193.980 0.000 194.360 0.380 ;
    END
  END din0[16]
  PIN din0[17]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 199.820 0.000 200.200 0.380 ;
    END
  END din0[17]
  PIN din0[18]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 205.660 0.000 206.040 0.380 ;
    END
  END din0[18]
  PIN din0[19]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 211.500 0.000 211.880 0.380 ;
    END
  END din0[19]
  PIN din0[20]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 217.340 0.000 217.720 0.380 ;
    END
  END din0[20]
  PIN din0[21]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 223.180 0.000 223.560 0.380 ;
    END
  END din0[21]
  PIN din0[22]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 229.020 0.000 229.400 0.380 ;
    END
  END din0[22]
  PIN din0[23]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 234.860 0.000 235.240 0.380 ;
    END
  END din0[23]
  PIN din0[24]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 240.700 0.000 241.080 0.380 ;
    END
  END din0[24]
  PIN din0[25]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 246.540 0.000 246.920 0.380 ;
    END
  END din0[25]
  PIN din0[26]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 252.380 0.000 252.760 0.380 ;
    END
  END din0[26]
  PIN din0[27]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 258.220 0.000 258.600 0.380 ;
    END
  END din0[27]
  PIN din0[28]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 264.060 0.000 264.440 0.380 ;
    END
  END din0[28]
  PIN din0[29]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 269.900 0.000 270.280 0.380 ;
    END
  END din0[29]
  PIN din0[30]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 275.740 0.000 276.120 0.380 ;
    END
  END din0[30]
  PIN din0[31]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 281.580 0.000 281.960 0.380 ;
    END
  END din0[31]
  PIN din0[32]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 287.420 0.000 287.800 0.380 ;
    END
  END din0[32]
  PIN addr0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 63.270 167.190 63.650 167.570 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 67.625 167.190 68.005 167.570 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 63.960 167.190 64.340 167.570 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 66.935 167.190 67.315 167.570 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 66.245 167.190 66.625 167.570 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 65.500 167.190 65.880 167.570 ;
    END
  END addr0[5]
  PIN csb0
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.830 0.380 23.210 ;
    END
  END csb0
  PIN web0
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.330 0.380 31.710 ;
    END
  END web0
  PIN clk0
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 31.100 0.000 31.480 0.380 ;
    END
  END clk0
  PIN wmask0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 77.180 0.000 77.560 0.380 ;
    END
  END wmask0[0]
  PIN wmask0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 83.020 0.000 83.400 0.380 ;
    END
  END wmask0[1]
  PIN wmask0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 88.860 0.000 89.240 0.380 ;
    END
  END wmask0[2]
  PIN wmask0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 94.700 0.000 95.080 0.380 ;
    END
  END wmask0[3]
  PIN spare_wen0
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 293.260 0.000 293.640 0.380 ;
    END
  END spare_wen0
  PIN dout0[0]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 131.225 0.000 131.605 0.380 ;
    END
  END dout0[0]
  PIN dout0[1]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 136.340 0.000 136.720 0.380 ;
    END
  END dout0[1]
  PIN dout0[2]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 137.490 0.000 137.870 0.380 ;
    END
  END dout0[2]
  PIN dout0[3]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 142.110 0.000 142.490 0.380 ;
    END
  END dout0[3]
  PIN dout0[4]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 143.870 0.000 144.250 0.380 ;
    END
  END dout0[4]
  PIN dout0[5]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 144.960 0.000 145.340 0.380 ;
    END
  END dout0[5]
  PIN dout0[6]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 147.950 0.000 148.330 0.380 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 149.960 0.000 150.340 0.380 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 153.870 0.000 154.250 0.380 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 156.340 0.000 156.720 0.380 ;
    END
  END dout0[9]
  PIN dout0[10]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 157.135 0.000 157.515 0.380 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 161.340 0.000 161.720 0.380 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 162.490 0.000 162.870 0.380 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 166.340 0.000 166.720 0.380 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 167.490 0.000 167.870 0.380 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 171.310 0.000 171.690 0.380 ;
    END
  END dout0[15]
  PIN dout0[16]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 173.870 0.000 174.250 0.380 ;
    END
  END dout0[16]
  PIN dout0[17]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 177.150 0.000 177.530 0.380 ;
    END
  END dout0[17]
  PIN dout0[18]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 178.870 0.000 179.250 0.380 ;
    END
  END dout0[18]
  PIN dout0[19]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 179.960 0.000 180.340 0.380 ;
    END
  END dout0[19]
  PIN dout0[20]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 182.990 0.000 183.370 0.380 ;
    END
  END dout0[20]
  PIN dout0[21]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 186.280 0.000 186.660 0.380 ;
    END
  END dout0[21]
  PIN dout0[22]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 188.870 0.000 189.250 0.380 ;
    END
  END dout0[22]
  PIN dout0[23]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 189.960 0.000 190.340 0.380 ;
    END
  END dout0[23]
  PIN dout0[24]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 194.670 0.000 195.050 0.380 ;
    END
  END dout0[24]
  PIN dout0[25]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 196.340 0.000 196.720 0.380 ;
    END
  END dout0[25]
  PIN dout0[26]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 197.490 0.000 197.870 0.380 ;
    END
  END dout0[26]
  PIN dout0[27]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 201.340 0.000 201.720 0.380 ;
    END
  END dout0[27]
  PIN dout0[28]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 202.490 0.000 202.870 0.380 ;
    END
  END dout0[28]
  PIN dout0[29]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 206.350 0.000 206.730 0.380 ;
    END
  END dout0[29]
  PIN dout0[30]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 207.490 0.000 207.870 0.380 ;
    END
  END dout0[30]
  PIN dout0[31]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 212.190 0.000 212.570 0.380 ;
    END
  END dout0[31]
  PIN dout0[32]
    DIRECTION OUTPUT ;
    PORT
      LAYER met4 ;
        RECT 215.035 0.000 215.415 0.380 ;
    END
  END dout0[32]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.740 167.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 0.000 310.680 1.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.940 0.000 310.680 167.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 165.830 310.680 167.570 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
        RECT 3.480 162.350 307.200 164.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.480 3.480 307.200 5.220 ;
    END
    PORT
      LAYER met4 ;
        RECT 305.460 3.480 307.200 164.090 ;
    END
    PORT
      LAYER met4 ;
        RECT 3.480 3.480 5.220 164.090 ;
    END
  END vssd1
  OBS
      LAYER met1 ;
        RECT 0.620 0.620 310.060 166.950 ;
      LAYER met2 ;
        RECT 0.620 0.620 310.060 166.950 ;
      LAYER met3 ;
        RECT 0.620 32.310 310.060 161.750 ;
        RECT 0.980 30.730 310.060 32.310 ;
        RECT 0.620 23.810 310.060 30.730 ;
        RECT 0.980 22.230 310.060 23.810 ;
        RECT 0.620 5.820 310.060 22.230 ;
      LAYER met4 ;
        RECT 5.830 166.590 62.670 166.950 ;
        RECT 68.605 166.590 304.880 166.950 ;
        RECT 5.830 164.690 304.880 166.590 ;
        RECT 5.830 5.820 304.860 164.690 ;
        RECT 5.830 0.980 49.730 5.820 ;
        RECT 5.830 0.620 30.500 0.980 ;
        RECT 32.080 0.620 49.730 0.980 ;
        RECT 70.790 0.980 295.450 5.820 ;
        RECT 70.790 0.620 76.580 0.980 ;
        RECT 78.160 0.620 82.420 0.980 ;
        RECT 84.000 0.620 88.260 0.980 ;
        RECT 89.840 0.620 94.100 0.980 ;
        RECT 95.680 0.620 99.940 0.980 ;
        RECT 101.520 0.620 105.780 0.980 ;
        RECT 107.360 0.620 111.620 0.980 ;
        RECT 113.200 0.620 117.460 0.980 ;
        RECT 119.040 0.620 123.300 0.980 ;
        RECT 124.880 0.620 129.140 0.980 ;
        RECT 132.205 0.620 134.980 0.980 ;
        RECT 138.470 0.620 140.820 0.980 ;
        RECT 143.090 0.620 143.270 0.980 ;
        RECT 145.940 0.620 146.660 0.980 ;
        RECT 148.930 0.620 149.360 0.980 ;
        RECT 150.940 0.620 152.500 0.980 ;
        RECT 154.850 0.620 155.740 0.980 ;
        RECT 158.115 0.620 158.340 0.980 ;
        RECT 159.920 0.620 160.740 0.980 ;
        RECT 163.470 0.620 164.180 0.980 ;
        RECT 168.470 0.620 170.020 0.980 ;
        RECT 172.290 0.620 173.270 0.980 ;
        RECT 174.850 0.620 175.860 0.980 ;
        RECT 178.130 0.620 178.270 0.980 ;
        RECT 180.940 0.620 181.700 0.980 ;
        RECT 183.970 0.620 185.680 0.980 ;
        RECT 187.260 0.620 187.540 0.980 ;
        RECT 190.940 0.620 193.380 0.980 ;
        RECT 195.650 0.620 195.740 0.980 ;
        RECT 198.470 0.620 199.220 0.980 ;
        RECT 203.470 0.620 205.060 0.980 ;
        RECT 208.470 0.620 210.900 0.980 ;
        RECT 213.170 0.620 214.435 0.980 ;
        RECT 216.015 0.620 216.740 0.980 ;
        RECT 218.320 0.620 222.580 0.980 ;
        RECT 224.160 0.620 228.420 0.980 ;
        RECT 230.000 0.620 234.260 0.980 ;
        RECT 235.840 0.620 240.100 0.980 ;
        RECT 241.680 0.620 245.940 0.980 ;
        RECT 247.520 0.620 251.780 0.980 ;
        RECT 253.360 0.620 257.620 0.980 ;
        RECT 259.200 0.620 263.460 0.980 ;
        RECT 265.040 0.620 269.300 0.980 ;
        RECT 270.880 0.620 275.140 0.980 ;
        RECT 276.720 0.620 280.980 0.980 ;
        RECT 282.560 0.620 286.820 0.980 ;
        RECT 288.400 0.620 292.660 0.980 ;
        RECT 294.240 0.620 295.450 0.980 ;
        RECT 304.860 0.620 304.880 2.880 ;
        RECT 34.010 0.610 49.730 0.620 ;
  END
END sky130_sram_256B_1rw_32x64
END LIBRARY

