module tt_um_openram_top (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire \dout[0] ;
 wire \dout[10] ;
 wire \dout[11] ;
 wire \dout[12] ;
 wire \dout[13] ;
 wire \dout[14] ;
 wire \dout[15] ;
 wire \dout[16] ;
 wire \dout[17] ;
 wire \dout[18] ;
 wire \dout[19] ;
 wire \dout[1] ;
 wire \dout[20] ;
 wire \dout[21] ;
 wire \dout[22] ;
 wire \dout[23] ;
 wire \dout[24] ;
 wire \dout[25] ;
 wire \dout[26] ;
 wire \dout[27] ;
 wire \dout[28] ;
 wire \dout[29] ;
 wire \dout[2] ;
 wire \dout[30] ;
 wire \dout[31] ;
 wire \dout[32] ;
 wire \dout[3] ;
 wire \dout[4] ;
 wire \dout[5] ;
 wire \dout[6] ;
 wire \dout[7] ;
 wire \dout[8] ;
 wire \dout[9] ;
 wire \scan_chain.scan_cells[0].scan_cell.data_out ;
 wire \scan_chain.scan_cells[0].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[10].scan_cell.data_out ;
 wire \scan_chain.scan_cells[10].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[10].scan_cell.scan_in ;
 wire \scan_chain.scan_cells[11].scan_cell.data_out ;
 wire \scan_chain.scan_cells[11].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[12].scan_cell.data_out ;
 wire \scan_chain.scan_cells[12].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[13].scan_cell.data_out ;
 wire \scan_chain.scan_cells[13].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[14].scan_cell.data_out ;
 wire \scan_chain.scan_cells[14].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[15].scan_cell.data_out ;
 wire \scan_chain.scan_cells[15].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[16].scan_cell.data_out ;
 wire \scan_chain.scan_cells[16].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[17].scan_cell.data_out ;
 wire \scan_chain.scan_cells[17].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[18].scan_cell.data_out ;
 wire \scan_chain.scan_cells[18].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[19].scan_cell.data_out ;
 wire \scan_chain.scan_cells[19].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[1].scan_cell.data_out ;
 wire \scan_chain.scan_cells[1].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[20].scan_cell.data_out ;
 wire \scan_chain.scan_cells[20].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[21].scan_cell.data_out ;
 wire \scan_chain.scan_cells[21].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[22].scan_cell.data_out ;
 wire \scan_chain.scan_cells[22].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[23].scan_cell.data_out ;
 wire \scan_chain.scan_cells[23].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[24].scan_cell.data_out ;
 wire \scan_chain.scan_cells[24].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[25].scan_cell.data_out ;
 wire \scan_chain.scan_cells[25].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[26].scan_cell.data_out ;
 wire \scan_chain.scan_cells[26].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[27].scan_cell.data_out ;
 wire \scan_chain.scan_cells[27].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[28].scan_cell.data_out ;
 wire \scan_chain.scan_cells[28].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[29].scan_cell.data_out ;
 wire \scan_chain.scan_cells[29].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[2].scan_cell.data_out ;
 wire \scan_chain.scan_cells[2].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[30].scan_cell.data_out ;
 wire \scan_chain.scan_cells[30].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[31].scan_cell.data_out ;
 wire \scan_chain.scan_cells[31].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[32].scan_cell.data_out ;
 wire \scan_chain.scan_cells[32].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[33].scan_cell.data_in ;
 wire \scan_chain.scan_cells[33].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[34].scan_cell.data_in ;
 wire \scan_chain.scan_cells[34].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[35].scan_cell.data_in ;
 wire \scan_chain.scan_cells[35].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[36].scan_cell.data_in ;
 wire \scan_chain.scan_cells[36].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[37].scan_cell.data_in ;
 wire \scan_chain.scan_cells[37].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[38].scan_cell.data_in ;
 wire \scan_chain.scan_cells[38].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[39].scan_cell.data_in ;
 wire \scan_chain.scan_cells[39].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[3].scan_cell.data_out ;
 wire \scan_chain.scan_cells[3].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[40].scan_cell.data_in ;
 wire \scan_chain.scan_cells[40].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[41].scan_cell.data_in ;
 wire \scan_chain.scan_cells[41].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[42].scan_cell.data_in ;
 wire \scan_chain.scan_cells[42].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[43].scan_cell.data_in ;
 wire \scan_chain.scan_cells[43].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[44].scan_cell.data_in ;
 wire \scan_chain.scan_cells[44].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[45].scan_cell.data_in ;
 wire \scan_chain.scan_cells[45].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[46].scan_cell.data_in ;
 wire \scan_chain.scan_cells[46].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[47].scan_cell.data_in ;
 wire \scan_chain.scan_cells[47].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[48].scan_cell.data_in ;
 wire \scan_chain.scan_cells[48].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[49].scan_cell.data_in ;
 wire \scan_chain.scan_cells[49].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[4].scan_cell.data_out ;
 wire \scan_chain.scan_cells[4].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[50].scan_cell.data_in ;
 wire \scan_chain.scan_cells[50].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[51].scan_cell.data_in ;
 wire \scan_chain.scan_cells[51].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[52].scan_cell.data_in ;
 wire \scan_chain.scan_cells[52].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[53].scan_cell.data_in ;
 wire \scan_chain.scan_cells[53].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[54].scan_cell.data_in ;
 wire \scan_chain.scan_cells[54].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[55].scan_cell.data_in ;
 wire \scan_chain.scan_cells[55].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[56].scan_cell.data_in ;
 wire \scan_chain.scan_cells[56].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[57].scan_cell.data_in ;
 wire \scan_chain.scan_cells[57].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[58].scan_cell.data_in ;
 wire \scan_chain.scan_cells[58].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[59].scan_cell.data_in ;
 wire \scan_chain.scan_cells[59].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[5].scan_cell.data_out ;
 wire \scan_chain.scan_cells[5].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[60].scan_cell.data_in ;
 wire \scan_chain.scan_cells[60].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[61].scan_cell.data_in ;
 wire \scan_chain.scan_cells[61].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[62].scan_cell.data_in ;
 wire \scan_chain.scan_cells[62].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[63].scan_cell.data_in ;
 wire \scan_chain.scan_cells[63].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[64].scan_cell.data_in ;
 wire \scan_chain.scan_cells[64].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[65].scan_cell.data_in ;
 wire \scan_chain.scan_cells[65].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[66].scan_cell.data_in ;
 wire \scan_chain.scan_cells[66].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[67].scan_cell.data_in ;
 wire \scan_chain.scan_cells[67].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[68].scan_cell.data_in ;
 wire \scan_chain.scan_cells[68].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[69].scan_cell.data_in ;
 wire \scan_chain.scan_cells[69].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[6].scan_cell.data_out ;
 wire \scan_chain.scan_cells[6].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[70].scan_cell.data_in ;
 wire \scan_chain.scan_cells[70].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[71].scan_cell.data_in ;
 wire \scan_chain.scan_cells[71].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[7].scan_cell.data_out ;
 wire \scan_chain.scan_cells[7].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[8].scan_cell.data_out ;
 wire \scan_chain.scan_cells[8].scan_cell.primary_ff ;
 wire \scan_chain.scan_cells[9].scan_cell.primary_ff ;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire [4:0] clknet_0_ui_in;
 wire [4:0] clknet_3_0__leaf_ui_in;
 wire [4:0] clknet_3_1__leaf_ui_in;
 wire [4:0] clknet_3_2__leaf_ui_in;
 wire [4:0] clknet_3_3__leaf_ui_in;
 wire [4:0] clknet_3_4__leaf_ui_in;
 wire [4:0] clknet_3_5__leaf_ui_in;
 wire [4:0] clknet_3_6__leaf_ui_in;
 wire [4:0] clknet_3_7__leaf_ui_in;

 sky130_sram_256B_1rw_32x64 SRAM (.csb0(ui_in[5]),
    .web0(ui_in[6]),
    .clk0(clknet_3_4__leaf_ui_in[3]),
    .spare_wen0(ui_in[7]),
    .addr0({\scan_chain.scan_cells[71].scan_cell.data_in ,
    \scan_chain.scan_cells[70].scan_cell.data_in ,
    \scan_chain.scan_cells[69].scan_cell.data_in ,
    \scan_chain.scan_cells[68].scan_cell.data_in ,
    \scan_chain.scan_cells[67].scan_cell.data_in ,
    \scan_chain.scan_cells[66].scan_cell.data_in }),
    .din0({\scan_chain.scan_cells[65].scan_cell.data_in ,
    \scan_chain.scan_cells[64].scan_cell.data_in ,
    \scan_chain.scan_cells[63].scan_cell.data_in ,
    \scan_chain.scan_cells[62].scan_cell.data_in ,
    \scan_chain.scan_cells[61].scan_cell.data_in ,
    \scan_chain.scan_cells[60].scan_cell.data_in ,
    \scan_chain.scan_cells[59].scan_cell.data_in ,
    \scan_chain.scan_cells[58].scan_cell.data_in ,
    \scan_chain.scan_cells[57].scan_cell.data_in ,
    \scan_chain.scan_cells[56].scan_cell.data_in ,
    \scan_chain.scan_cells[55].scan_cell.data_in ,
    \scan_chain.scan_cells[54].scan_cell.data_in ,
    \scan_chain.scan_cells[53].scan_cell.data_in ,
    \scan_chain.scan_cells[52].scan_cell.data_in ,
    \scan_chain.scan_cells[51].scan_cell.data_in ,
    \scan_chain.scan_cells[50].scan_cell.data_in ,
    \scan_chain.scan_cells[49].scan_cell.data_in ,
    \scan_chain.scan_cells[48].scan_cell.data_in ,
    \scan_chain.scan_cells[47].scan_cell.data_in ,
    \scan_chain.scan_cells[46].scan_cell.data_in ,
    \scan_chain.scan_cells[45].scan_cell.data_in ,
    \scan_chain.scan_cells[44].scan_cell.data_in ,
    \scan_chain.scan_cells[43].scan_cell.data_in ,
    \scan_chain.scan_cells[42].scan_cell.data_in ,
    \scan_chain.scan_cells[41].scan_cell.data_in ,
    \scan_chain.scan_cells[40].scan_cell.data_in ,
    \scan_chain.scan_cells[39].scan_cell.data_in ,
    \scan_chain.scan_cells[38].scan_cell.data_in ,
    \scan_chain.scan_cells[37].scan_cell.data_in ,
    \scan_chain.scan_cells[36].scan_cell.data_in ,
    \scan_chain.scan_cells[35].scan_cell.data_in ,
    \scan_chain.scan_cells[34].scan_cell.data_in ,
    \scan_chain.scan_cells[33].scan_cell.data_in }),
    .dout0({\dout[32] ,
    \dout[31] ,
    \dout[30] ,
    \dout[29] ,
    \dout[28] ,
    \dout[27] ,
    \dout[26] ,
    \dout[25] ,
    \dout[24] ,
    \dout[23] ,
    \dout[22] ,
    \dout[21] ,
    \dout[20] ,
    \dout[19] ,
    \dout[18] ,
    \dout[17] ,
    \dout[16] ,
    \dout[15] ,
    \dout[14] ,
    \dout[13] ,
    \dout[12] ,
    \dout[11] ,
    \dout[10] ,
    \dout[9] ,
    \dout[8] ,
    \dout[7] ,
    \dout[6] ,
    \dout[5] ,
    \dout[4] ,
    \dout[3] ,
    \dout[2] ,
    \dout[1] ,
    \dout[0] }),
    .wmask0({uio_in[3],
    uio_in[2],
    uio_in[1],
    uio_in[0]}));
 sky130_fd_sc_hd__mux2_1 _250_ (.A0(\scan_chain.scan_cells[10].scan_cell.scan_in ),
    .A1(\scan_chain.scan_cells[8].scan_cell.data_out ),
    .S(net12),
    .X(_144_));
 sky130_fd_sc_hd__mux2_1 _251_ (.A0(\scan_chain.scan_cells[9].scan_cell.primary_ff ),
    .A1(_144_),
    .S(net27),
    .X(_026_));
 sky130_fd_sc_hd__nand2_2 _252_ (.A(net20),
    .B(net34),
    .Y(_145_));
 sky130_fd_sc_hd__mux2_1 _253_ (.A0(\scan_chain.scan_cells[71].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[71].scan_cell.data_in ),
    .S(net5),
    .X(_027_));
 sky130_fd_sc_hd__mux2_1 _254_ (.A0(\scan_chain.scan_cells[70].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[69].scan_cell.data_in ),
    .S(net9),
    .X(_146_));
 sky130_fd_sc_hd__mux2_1 _255_ (.A0(\scan_chain.scan_cells[70].scan_cell.primary_ff ),
    .A1(_146_),
    .S(net25),
    .X(_028_));
 sky130_fd_sc_hd__mux2_1 _256_ (.A0(\scan_chain.scan_cells[70].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[70].scan_cell.data_in ),
    .S(net5),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _257_ (.A0(\scan_chain.scan_cells[6].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[5].scan_cell.data_out ),
    .S(net10),
    .X(_147_));
 sky130_fd_sc_hd__mux2_1 _258_ (.A0(\scan_chain.scan_cells[6].scan_cell.primary_ff ),
    .A1(_147_),
    .S(net23),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _259_ (.A0(\scan_chain.scan_cells[69].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[69].scan_cell.data_in ),
    .S(net5),
    .X(_031_));
 sky130_fd_sc_hd__mux2_1 _260_ (.A0(\scan_chain.scan_cells[68].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[67].scan_cell.data_in ),
    .S(net9),
    .X(_148_));
 sky130_fd_sc_hd__mux2_1 _261_ (.A0(\scan_chain.scan_cells[68].scan_cell.primary_ff ),
    .A1(_148_),
    .S(net25),
    .X(_032_));
 sky130_fd_sc_hd__mux2_1 _262_ (.A0(\scan_chain.scan_cells[68].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[68].scan_cell.data_in ),
    .S(net5),
    .X(_033_));
 sky130_fd_sc_hd__mux2_1 _263_ (.A0(\scan_chain.scan_cells[67].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[66].scan_cell.data_in ),
    .S(net9),
    .X(_149_));
 sky130_fd_sc_hd__mux2_1 _264_ (.A0(\scan_chain.scan_cells[67].scan_cell.primary_ff ),
    .A1(_149_),
    .S(net25),
    .X(_034_));
 sky130_fd_sc_hd__mux2_1 _265_ (.A0(\scan_chain.scan_cells[67].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[67].scan_cell.data_in ),
    .S(net5),
    .X(_035_));
 sky130_fd_sc_hd__mux2_1 _266_ (.A0(\scan_chain.scan_cells[66].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[65].scan_cell.data_in ),
    .S(net9),
    .X(_150_));
 sky130_fd_sc_hd__mux2_1 _267_ (.A0(\scan_chain.scan_cells[66].scan_cell.primary_ff ),
    .A1(_150_),
    .S(net25),
    .X(_036_));
 sky130_fd_sc_hd__mux2_1 _268_ (.A0(\scan_chain.scan_cells[66].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[66].scan_cell.data_in ),
    .S(net5),
    .X(_037_));
 sky130_fd_sc_hd__mux2_1 _269_ (.A0(\scan_chain.scan_cells[65].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[64].scan_cell.data_in ),
    .S(net20),
    .X(_151_));
 sky130_fd_sc_hd__mux2_1 _270_ (.A0(\scan_chain.scan_cells[65].scan_cell.primary_ff ),
    .A1(_151_),
    .S(net34),
    .X(_038_));
 sky130_fd_sc_hd__mux2_1 _271_ (.A0(\scan_chain.scan_cells[65].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[65].scan_cell.data_in ),
    .S(net7),
    .X(_039_));
 sky130_fd_sc_hd__mux2_1 _272_ (.A0(\scan_chain.scan_cells[64].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[63].scan_cell.data_in ),
    .S(net20),
    .X(_152_));
 sky130_fd_sc_hd__mux2_1 _273_ (.A0(\scan_chain.scan_cells[64].scan_cell.primary_ff ),
    .A1(_152_),
    .S(net34),
    .X(_040_));
 sky130_fd_sc_hd__mux2_1 _274_ (.A0(\scan_chain.scan_cells[64].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[64].scan_cell.data_in ),
    .S(net8),
    .X(_041_));
 sky130_fd_sc_hd__mux2_1 _275_ (.A0(\scan_chain.scan_cells[63].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[62].scan_cell.data_in ),
    .S(net20),
    .X(_153_));
 sky130_fd_sc_hd__mux2_1 _276_ (.A0(\scan_chain.scan_cells[63].scan_cell.primary_ff ),
    .A1(_153_),
    .S(net34),
    .X(_042_));
 sky130_fd_sc_hd__mux2_1 _277_ (.A0(\scan_chain.scan_cells[63].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[63].scan_cell.data_in ),
    .S(net7),
    .X(_043_));
 sky130_fd_sc_hd__mux2_1 _278_ (.A0(\scan_chain.scan_cells[62].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[61].scan_cell.data_in ),
    .S(net21),
    .X(_154_));
 sky130_fd_sc_hd__mux2_1 _279_ (.A0(\scan_chain.scan_cells[62].scan_cell.primary_ff ),
    .A1(_154_),
    .S(net34),
    .X(_044_));
 sky130_fd_sc_hd__mux2_1 _280_ (.A0(\scan_chain.scan_cells[62].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[62].scan_cell.data_in ),
    .S(net7),
    .X(_045_));
 sky130_fd_sc_hd__mux2_1 _281_ (.A0(\scan_chain.scan_cells[61].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[60].scan_cell.data_in ),
    .S(net21),
    .X(_155_));
 sky130_fd_sc_hd__mux2_1 _282_ (.A0(\scan_chain.scan_cells[61].scan_cell.primary_ff ),
    .A1(_155_),
    .S(net34),
    .X(_046_));
 sky130_fd_sc_hd__mux2_1 _283_ (.A0(\scan_chain.scan_cells[61].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[61].scan_cell.data_in ),
    .S(net7),
    .X(_047_));
 sky130_fd_sc_hd__mux2_1 _284_ (.A0(\scan_chain.scan_cells[60].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[59].scan_cell.data_in ),
    .S(net21),
    .X(_156_));
 sky130_fd_sc_hd__mux2_1 _285_ (.A0(\scan_chain.scan_cells[60].scan_cell.primary_ff ),
    .A1(_156_),
    .S(net34),
    .X(_048_));
 sky130_fd_sc_hd__mux2_1 _286_ (.A0(\scan_chain.scan_cells[60].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[60].scan_cell.data_in ),
    .S(net7),
    .X(_049_));
 sky130_fd_sc_hd__mux2_1 _287_ (.A0(\scan_chain.scan_cells[5].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[4].scan_cell.data_out ),
    .S(net10),
    .X(_157_));
 sky130_fd_sc_hd__mux2_1 _288_ (.A0(\scan_chain.scan_cells[5].scan_cell.primary_ff ),
    .A1(_157_),
    .S(net23),
    .X(_050_));
 sky130_fd_sc_hd__mux2_1 _289_ (.A0(\scan_chain.scan_cells[59].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[59].scan_cell.data_in ),
    .S(net7),
    .X(_051_));
 sky130_fd_sc_hd__mux2_1 _290_ (.A0(\scan_chain.scan_cells[58].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[57].scan_cell.data_in ),
    .S(net18),
    .X(_158_));
 sky130_fd_sc_hd__mux2_1 _291_ (.A0(\scan_chain.scan_cells[58].scan_cell.primary_ff ),
    .A1(_158_),
    .S(net33),
    .X(_052_));
 sky130_fd_sc_hd__mux2_1 _292_ (.A0(\scan_chain.scan_cells[58].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[58].scan_cell.data_in ),
    .S(net7),
    .X(_053_));
 sky130_fd_sc_hd__mux2_1 _293_ (.A0(\scan_chain.scan_cells[57].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[56].scan_cell.data_in ),
    .S(net18),
    .X(_159_));
 sky130_fd_sc_hd__mux2_1 _294_ (.A0(\scan_chain.scan_cells[57].scan_cell.primary_ff ),
    .A1(_159_),
    .S(net33),
    .X(_054_));
 sky130_fd_sc_hd__mux2_1 _295_ (.A0(\scan_chain.scan_cells[57].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[57].scan_cell.data_in ),
    .S(net7),
    .X(_055_));
 sky130_fd_sc_hd__mux2_1 _296_ (.A0(\scan_chain.scan_cells[56].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[55].scan_cell.data_in ),
    .S(net18),
    .X(_160_));
 sky130_fd_sc_hd__mux2_1 _297_ (.A0(\scan_chain.scan_cells[56].scan_cell.primary_ff ),
    .A1(_160_),
    .S(net33),
    .X(_056_));
 sky130_fd_sc_hd__mux2_1 _298_ (.A0(\scan_chain.scan_cells[56].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[56].scan_cell.data_in ),
    .S(net7),
    .X(_057_));
 sky130_fd_sc_hd__mux2_1 _299_ (.A0(\scan_chain.scan_cells[55].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[54].scan_cell.data_in ),
    .S(net18),
    .X(_161_));
 sky130_fd_sc_hd__mux2_1 _300_ (.A0(\scan_chain.scan_cells[55].scan_cell.primary_ff ),
    .A1(_161_),
    .S(net33),
    .X(_058_));
 sky130_fd_sc_hd__mux2_1 _301_ (.A0(\scan_chain.scan_cells[55].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[55].scan_cell.data_in ),
    .S(net8),
    .X(_059_));
 sky130_fd_sc_hd__mux2_1 _302_ (.A0(\scan_chain.scan_cells[54].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[53].scan_cell.data_in ),
    .S(net18),
    .X(_162_));
 sky130_fd_sc_hd__mux2_1 _303_ (.A0(\scan_chain.scan_cells[54].scan_cell.primary_ff ),
    .A1(_162_),
    .S(net33),
    .X(_060_));
 sky130_fd_sc_hd__mux2_1 _304_ (.A0(\scan_chain.scan_cells[54].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[54].scan_cell.data_in ),
    .S(net7),
    .X(_061_));
 sky130_fd_sc_hd__mux2_1 _305_ (.A0(\scan_chain.scan_cells[53].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[52].scan_cell.data_in ),
    .S(net18),
    .X(_163_));
 sky130_fd_sc_hd__mux2_1 _306_ (.A0(\scan_chain.scan_cells[53].scan_cell.primary_ff ),
    .A1(_163_),
    .S(net33),
    .X(_062_));
 sky130_fd_sc_hd__mux2_1 _307_ (.A0(\scan_chain.scan_cells[53].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[53].scan_cell.data_in ),
    .S(net8),
    .X(_063_));
 sky130_fd_sc_hd__mux2_1 _308_ (.A0(\scan_chain.scan_cells[52].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[51].scan_cell.data_in ),
    .S(net17),
    .X(_164_));
 sky130_fd_sc_hd__mux2_1 _309_ (.A0(\scan_chain.scan_cells[52].scan_cell.primary_ff ),
    .A1(_164_),
    .S(net32),
    .X(_064_));
 sky130_fd_sc_hd__mux2_1 _310_ (.A0(\scan_chain.scan_cells[52].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[52].scan_cell.data_in ),
    .S(net8),
    .X(_065_));
 sky130_fd_sc_hd__mux2_1 _311_ (.A0(\scan_chain.scan_cells[51].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[50].scan_cell.data_in ),
    .S(net17),
    .X(_165_));
 sky130_fd_sc_hd__mux2_1 _312_ (.A0(\scan_chain.scan_cells[51].scan_cell.primary_ff ),
    .A1(_165_),
    .S(net31),
    .X(_066_));
 sky130_fd_sc_hd__mux2_1 _313_ (.A0(\scan_chain.scan_cells[51].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[51].scan_cell.data_in ),
    .S(net8),
    .X(_067_));
 sky130_fd_sc_hd__mux2_1 _314_ (.A0(\scan_chain.scan_cells[50].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[49].scan_cell.data_in ),
    .S(net17),
    .X(_166_));
 sky130_fd_sc_hd__mux2_1 _315_ (.A0(\scan_chain.scan_cells[50].scan_cell.primary_ff ),
    .A1(_166_),
    .S(net31),
    .X(_068_));
 sky130_fd_sc_hd__mux2_1 _316_ (.A0(\scan_chain.scan_cells[50].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[50].scan_cell.data_in ),
    .S(net8),
    .X(_069_));
 sky130_fd_sc_hd__mux2_1 _317_ (.A0(\scan_chain.scan_cells[4].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[3].scan_cell.data_out ),
    .S(net9),
    .X(_167_));
 sky130_fd_sc_hd__mux2_1 _318_ (.A0(\scan_chain.scan_cells[4].scan_cell.primary_ff ),
    .A1(_167_),
    .S(net23),
    .X(_070_));
 sky130_fd_sc_hd__mux2_1 _319_ (.A0(\scan_chain.scan_cells[49].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[49].scan_cell.data_in ),
    .S(net8),
    .X(_071_));
 sky130_fd_sc_hd__mux2_1 _320_ (.A0(\scan_chain.scan_cells[48].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[47].scan_cell.data_in ),
    .S(net13),
    .X(_168_));
 sky130_fd_sc_hd__mux2_1 _321_ (.A0(\scan_chain.scan_cells[48].scan_cell.primary_ff ),
    .A1(_168_),
    .S(net31),
    .X(_072_));
 sky130_fd_sc_hd__mux2_1 _322_ (.A0(\scan_chain.scan_cells[48].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[48].scan_cell.data_in ),
    .S(net8),
    .X(_073_));
 sky130_fd_sc_hd__mux2_1 _323_ (.A0(\scan_chain.scan_cells[47].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[46].scan_cell.data_in ),
    .S(net13),
    .X(_169_));
 sky130_fd_sc_hd__mux2_1 _324_ (.A0(\scan_chain.scan_cells[47].scan_cell.primary_ff ),
    .A1(_169_),
    .S(net28),
    .X(_074_));
 sky130_fd_sc_hd__mux2_1 _325_ (.A0(\scan_chain.scan_cells[47].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[47].scan_cell.data_in ),
    .S(net8),
    .X(_075_));
 sky130_fd_sc_hd__mux2_1 _326_ (.A0(\scan_chain.scan_cells[46].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[45].scan_cell.data_in ),
    .S(net13),
    .X(_170_));
 sky130_fd_sc_hd__mux2_1 _327_ (.A0(\scan_chain.scan_cells[46].scan_cell.primary_ff ),
    .A1(_170_),
    .S(net28),
    .X(_076_));
 sky130_fd_sc_hd__mux2_1 _328_ (.A0(\scan_chain.scan_cells[46].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[46].scan_cell.data_in ),
    .S(net6),
    .X(_077_));
 sky130_fd_sc_hd__mux2_1 _329_ (.A0(\scan_chain.scan_cells[45].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[44].scan_cell.data_in ),
    .S(net12),
    .X(_171_));
 sky130_fd_sc_hd__mux2_1 _330_ (.A0(\scan_chain.scan_cells[45].scan_cell.primary_ff ),
    .A1(_171_),
    .S(net27),
    .X(_078_));
 sky130_fd_sc_hd__mux2_1 _331_ (.A0(\scan_chain.scan_cells[45].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[45].scan_cell.data_in ),
    .S(net6),
    .X(_079_));
 sky130_fd_sc_hd__mux2_1 _332_ (.A0(\scan_chain.scan_cells[44].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[43].scan_cell.data_in ),
    .S(net12),
    .X(_172_));
 sky130_fd_sc_hd__mux2_1 _333_ (.A0(\scan_chain.scan_cells[44].scan_cell.primary_ff ),
    .A1(_172_),
    .S(net27),
    .X(_080_));
 sky130_fd_sc_hd__mux2_1 _334_ (.A0(\scan_chain.scan_cells[44].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[44].scan_cell.data_in ),
    .S(net6),
    .X(_081_));
 sky130_fd_sc_hd__mux2_1 _335_ (.A0(\scan_chain.scan_cells[43].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[42].scan_cell.data_in ),
    .S(net12),
    .X(_173_));
 sky130_fd_sc_hd__mux2_1 _336_ (.A0(\scan_chain.scan_cells[43].scan_cell.primary_ff ),
    .A1(_173_),
    .S(net27),
    .X(_082_));
 sky130_fd_sc_hd__mux2_1 _337_ (.A0(\scan_chain.scan_cells[43].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[43].scan_cell.data_in ),
    .S(net6),
    .X(_083_));
 sky130_fd_sc_hd__mux2_1 _338_ (.A0(\scan_chain.scan_cells[42].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[41].scan_cell.data_in ),
    .S(net12),
    .X(_174_));
 sky130_fd_sc_hd__mux2_1 _339_ (.A0(\scan_chain.scan_cells[42].scan_cell.primary_ff ),
    .A1(_174_),
    .S(net27),
    .X(_084_));
 sky130_fd_sc_hd__mux2_1 _340_ (.A0(\scan_chain.scan_cells[42].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[42].scan_cell.data_in ),
    .S(net6),
    .X(_085_));
 sky130_fd_sc_hd__mux2_1 _341_ (.A0(\scan_chain.scan_cells[41].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[40].scan_cell.data_in ),
    .S(net12),
    .X(_175_));
 sky130_fd_sc_hd__mux2_1 _342_ (.A0(\scan_chain.scan_cells[41].scan_cell.primary_ff ),
    .A1(_175_),
    .S(net27),
    .X(_086_));
 sky130_fd_sc_hd__mux2_1 _343_ (.A0(\scan_chain.scan_cells[41].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[41].scan_cell.data_in ),
    .S(_145_),
    .X(_087_));
 sky130_fd_sc_hd__mux2_1 _344_ (.A0(\scan_chain.scan_cells[40].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[39].scan_cell.data_in ),
    .S(net12),
    .X(_176_));
 sky130_fd_sc_hd__mux2_1 _345_ (.A0(\scan_chain.scan_cells[40].scan_cell.primary_ff ),
    .A1(_176_),
    .S(net27),
    .X(_088_));
 sky130_fd_sc_hd__mux2_1 _346_ (.A0(\scan_chain.scan_cells[40].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[40].scan_cell.data_in ),
    .S(net6),
    .X(_089_));
 sky130_fd_sc_hd__mux2_1 _347_ (.A0(\scan_chain.scan_cells[3].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[2].scan_cell.data_out ),
    .S(net9),
    .X(_177_));
 sky130_fd_sc_hd__mux2_1 _348_ (.A0(\scan_chain.scan_cells[3].scan_cell.primary_ff ),
    .A1(_177_),
    .S(net23),
    .X(_090_));
 sky130_fd_sc_hd__mux2_1 _349_ (.A0(\scan_chain.scan_cells[39].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[39].scan_cell.data_in ),
    .S(net6),
    .X(_091_));
 sky130_fd_sc_hd__mux2_1 _350_ (.A0(\scan_chain.scan_cells[38].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[37].scan_cell.data_in ),
    .S(net11),
    .X(_178_));
 sky130_fd_sc_hd__mux2_1 _351_ (.A0(\scan_chain.scan_cells[38].scan_cell.primary_ff ),
    .A1(_178_),
    .S(net26),
    .X(_092_));
 sky130_fd_sc_hd__mux2_1 _352_ (.A0(\scan_chain.scan_cells[38].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[38].scan_cell.data_in ),
    .S(net6),
    .X(_093_));
 sky130_fd_sc_hd__mux2_1 _353_ (.A0(\scan_chain.scan_cells[37].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[36].scan_cell.data_in ),
    .S(net11),
    .X(_179_));
 sky130_fd_sc_hd__mux2_1 _354_ (.A0(\scan_chain.scan_cells[37].scan_cell.primary_ff ),
    .A1(_179_),
    .S(net26),
    .X(_094_));
 sky130_fd_sc_hd__mux2_1 _355_ (.A0(\scan_chain.scan_cells[37].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[37].scan_cell.data_in ),
    .S(net5),
    .X(_095_));
 sky130_fd_sc_hd__mux2_1 _356_ (.A0(\scan_chain.scan_cells[36].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[35].scan_cell.data_in ),
    .S(net9),
    .X(_180_));
 sky130_fd_sc_hd__mux2_1 _357_ (.A0(\scan_chain.scan_cells[36].scan_cell.primary_ff ),
    .A1(_180_),
    .S(net25),
    .X(_096_));
 sky130_fd_sc_hd__mux2_1 _358_ (.A0(\scan_chain.scan_cells[36].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[36].scan_cell.data_in ),
    .S(net6),
    .X(_097_));
 sky130_fd_sc_hd__mux2_1 _359_ (.A0(\scan_chain.scan_cells[35].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[34].scan_cell.data_in ),
    .S(net9),
    .X(_181_));
 sky130_fd_sc_hd__mux2_1 _360_ (.A0(\scan_chain.scan_cells[35].scan_cell.primary_ff ),
    .A1(_181_),
    .S(net25),
    .X(_098_));
 sky130_fd_sc_hd__mux2_1 _361_ (.A0(\scan_chain.scan_cells[35].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[35].scan_cell.data_in ),
    .S(net5),
    .X(_099_));
 sky130_fd_sc_hd__mux2_1 _362_ (.A0(\scan_chain.scan_cells[34].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[33].scan_cell.data_in ),
    .S(net9),
    .X(_182_));
 sky130_fd_sc_hd__mux2_1 _363_ (.A0(\scan_chain.scan_cells[34].scan_cell.primary_ff ),
    .A1(_182_),
    .S(net25),
    .X(_100_));
 sky130_fd_sc_hd__mux2_1 _364_ (.A0(\scan_chain.scan_cells[34].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[34].scan_cell.data_in ),
    .S(net5),
    .X(_101_));
 sky130_fd_sc_hd__mux2_1 _365_ (.A0(\scan_chain.scan_cells[33].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[32].scan_cell.data_out ),
    .S(net9),
    .X(_183_));
 sky130_fd_sc_hd__mux2_1 _366_ (.A0(\scan_chain.scan_cells[33].scan_cell.primary_ff ),
    .A1(_183_),
    .S(net25),
    .X(_102_));
 sky130_fd_sc_hd__mux2_1 _367_ (.A0(\scan_chain.scan_cells[33].scan_cell.primary_ff ),
    .A1(\scan_chain.scan_cells[33].scan_cell.data_in ),
    .S(net5),
    .X(_103_));
 sky130_fd_sc_hd__mux2_1 _368_ (.A0(\scan_chain.scan_cells[32].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[31].scan_cell.data_out ),
    .S(net17),
    .X(_184_));
 sky130_fd_sc_hd__mux2_1 _369_ (.A0(\scan_chain.scan_cells[32].scan_cell.primary_ff ),
    .A1(_184_),
    .S(net31),
    .X(_104_));
 sky130_fd_sc_hd__mux2_1 _370_ (.A0(\dout[32] ),
    .A1(\scan_chain.scan_cells[32].scan_cell.primary_ff ),
    .S(net17),
    .X(_185_));
 sky130_fd_sc_hd__mux2_1 _371_ (.A0(\scan_chain.scan_cells[32].scan_cell.data_out ),
    .A1(_185_),
    .S(net32),
    .X(_105_));
 sky130_fd_sc_hd__mux2_1 _372_ (.A0(\scan_chain.scan_cells[31].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[30].scan_cell.data_out ),
    .S(net17),
    .X(_186_));
 sky130_fd_sc_hd__mux2_1 _373_ (.A0(\scan_chain.scan_cells[31].scan_cell.primary_ff ),
    .A1(_186_),
    .S(net32),
    .X(_106_));
 sky130_fd_sc_hd__mux2_1 _374_ (.A0(\dout[31] ),
    .A1(\scan_chain.scan_cells[31].scan_cell.primary_ff ),
    .S(net17),
    .X(_187_));
 sky130_fd_sc_hd__mux2_1 _375_ (.A0(\scan_chain.scan_cells[31].scan_cell.data_out ),
    .A1(_187_),
    .S(net32),
    .X(_107_));
 sky130_fd_sc_hd__mux2_1 _376_ (.A0(\scan_chain.scan_cells[30].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[29].scan_cell.data_out ),
    .S(net18),
    .X(_188_));
 sky130_fd_sc_hd__mux2_1 _377_ (.A0(\scan_chain.scan_cells[30].scan_cell.primary_ff ),
    .A1(_188_),
    .S(net33),
    .X(_108_));
 sky130_fd_sc_hd__mux2_1 _378_ (.A0(\dout[30] ),
    .A1(\scan_chain.scan_cells[30].scan_cell.primary_ff ),
    .S(net17),
    .X(_189_));
 sky130_fd_sc_hd__mux2_1 _379_ (.A0(\scan_chain.scan_cells[30].scan_cell.data_out ),
    .A1(_189_),
    .S(net36),
    .X(_109_));
 sky130_fd_sc_hd__mux2_1 _380_ (.A0(\scan_chain.scan_cells[2].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[1].scan_cell.data_out ),
    .S(net10),
    .X(_190_));
 sky130_fd_sc_hd__mux2_1 _381_ (.A0(\scan_chain.scan_cells[2].scan_cell.primary_ff ),
    .A1(_190_),
    .S(net23),
    .X(_110_));
 sky130_fd_sc_hd__mux2_1 _382_ (.A0(\dout[29] ),
    .A1(\scan_chain.scan_cells[29].scan_cell.primary_ff ),
    .S(net18),
    .X(_191_));
 sky130_fd_sc_hd__mux2_1 _383_ (.A0(\scan_chain.scan_cells[29].scan_cell.data_out ),
    .A1(_191_),
    .S(net33),
    .X(_111_));
 sky130_fd_sc_hd__mux2_1 _384_ (.A0(\scan_chain.scan_cells[28].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[27].scan_cell.data_out ),
    .S(net21),
    .X(_192_));
 sky130_fd_sc_hd__mux2_1 _385_ (.A0(\scan_chain.scan_cells[28].scan_cell.primary_ff ),
    .A1(_192_),
    .S(net34),
    .X(_112_));
 sky130_fd_sc_hd__mux2_1 _386_ (.A0(\dout[28] ),
    .A1(\scan_chain.scan_cells[28].scan_cell.primary_ff ),
    .S(net18),
    .X(_193_));
 sky130_fd_sc_hd__mux2_1 _387_ (.A0(\scan_chain.scan_cells[28].scan_cell.data_out ),
    .A1(_193_),
    .S(net33),
    .X(_113_));
 sky130_fd_sc_hd__mux2_1 _388_ (.A0(\scan_chain.scan_cells[27].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[26].scan_cell.data_out ),
    .S(net20),
    .X(_194_));
 sky130_fd_sc_hd__mux2_1 _389_ (.A0(\scan_chain.scan_cells[27].scan_cell.primary_ff ),
    .A1(_194_),
    .S(net35),
    .X(_114_));
 sky130_fd_sc_hd__mux2_1 _390_ (.A0(\dout[27] ),
    .A1(\scan_chain.scan_cells[27].scan_cell.primary_ff ),
    .S(net20),
    .X(_195_));
 sky130_fd_sc_hd__mux2_1 _391_ (.A0(\scan_chain.scan_cells[27].scan_cell.data_out ),
    .A1(_195_),
    .S(net34),
    .X(_115_));
 sky130_fd_sc_hd__mux2_1 _392_ (.A0(\scan_chain.scan_cells[26].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[25].scan_cell.data_out ),
    .S(net16),
    .X(_196_));
 sky130_fd_sc_hd__mux2_1 _393_ (.A0(\scan_chain.scan_cells[26].scan_cell.primary_ff ),
    .A1(_196_),
    .S(net30),
    .X(_116_));
 sky130_fd_sc_hd__mux2_1 _394_ (.A0(\dout[26] ),
    .A1(\scan_chain.scan_cells[26].scan_cell.primary_ff ),
    .S(net16),
    .X(_197_));
 sky130_fd_sc_hd__mux2_1 _395_ (.A0(\scan_chain.scan_cells[26].scan_cell.data_out ),
    .A1(_197_),
    .S(net30),
    .X(_117_));
 sky130_fd_sc_hd__mux2_1 _396_ (.A0(\scan_chain.scan_cells[25].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[24].scan_cell.data_out ),
    .S(net16),
    .X(_198_));
 sky130_fd_sc_hd__mux2_1 _397_ (.A0(\scan_chain.scan_cells[25].scan_cell.primary_ff ),
    .A1(_198_),
    .S(net30),
    .X(_118_));
 sky130_fd_sc_hd__mux2_1 _398_ (.A0(\dout[25] ),
    .A1(\scan_chain.scan_cells[25].scan_cell.primary_ff ),
    .S(net16),
    .X(_199_));
 sky130_fd_sc_hd__mux2_1 _399_ (.A0(\scan_chain.scan_cells[25].scan_cell.data_out ),
    .A1(_199_),
    .S(net30),
    .X(_119_));
 sky130_fd_sc_hd__mux2_1 _400_ (.A0(\scan_chain.scan_cells[24].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[23].scan_cell.data_out ),
    .S(net16),
    .X(_200_));
 sky130_fd_sc_hd__mux2_1 _401_ (.A0(\scan_chain.scan_cells[24].scan_cell.primary_ff ),
    .A1(_200_),
    .S(net30),
    .X(_120_));
 sky130_fd_sc_hd__mux2_1 _402_ (.A0(\dout[24] ),
    .A1(\scan_chain.scan_cells[24].scan_cell.primary_ff ),
    .S(net16),
    .X(_201_));
 sky130_fd_sc_hd__mux2_1 _403_ (.A0(\scan_chain.scan_cells[24].scan_cell.data_out ),
    .A1(_201_),
    .S(net30),
    .X(_121_));
 sky130_fd_sc_hd__mux2_1 _404_ (.A0(\scan_chain.scan_cells[23].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[22].scan_cell.data_out ),
    .S(net22),
    .X(_202_));
 sky130_fd_sc_hd__mux2_1 _405_ (.A0(\scan_chain.scan_cells[23].scan_cell.primary_ff ),
    .A1(_202_),
    .S(net30),
    .X(_122_));
 sky130_fd_sc_hd__mux2_1 _406_ (.A0(\dout[23] ),
    .A1(\scan_chain.scan_cells[23].scan_cell.primary_ff ),
    .S(net22),
    .X(_203_));
 sky130_fd_sc_hd__mux2_1 _407_ (.A0(\scan_chain.scan_cells[23].scan_cell.data_out ),
    .A1(_203_),
    .S(net37),
    .X(_123_));
 sky130_fd_sc_hd__mux2_1 _408_ (.A0(\scan_chain.scan_cells[22].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[21].scan_cell.data_out ),
    .S(net20),
    .X(_204_));
 sky130_fd_sc_hd__mux2_1 _409_ (.A0(\scan_chain.scan_cells[22].scan_cell.primary_ff ),
    .A1(_204_),
    .S(net35),
    .X(_124_));
 sky130_fd_sc_hd__mux2_1 _410_ (.A0(\dout[22] ),
    .A1(\scan_chain.scan_cells[22].scan_cell.primary_ff ),
    .S(net20),
    .X(_205_));
 sky130_fd_sc_hd__mux2_1 _411_ (.A0(\scan_chain.scan_cells[22].scan_cell.data_out ),
    .A1(_205_),
    .S(net35),
    .X(_125_));
 sky130_fd_sc_hd__mux2_1 _412_ (.A0(\scan_chain.scan_cells[21].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[20].scan_cell.data_out ),
    .S(net20),
    .X(_206_));
 sky130_fd_sc_hd__mux2_1 _413_ (.A0(\scan_chain.scan_cells[21].scan_cell.primary_ff ),
    .A1(_206_),
    .S(net35),
    .X(_126_));
 sky130_fd_sc_hd__mux2_1 _414_ (.A0(\dout[21] ),
    .A1(\scan_chain.scan_cells[21].scan_cell.primary_ff ),
    .S(net20),
    .X(_207_));
 sky130_fd_sc_hd__mux2_1 _415_ (.A0(\scan_chain.scan_cells[21].scan_cell.data_out ),
    .A1(_207_),
    .S(net35),
    .X(_127_));
 sky130_fd_sc_hd__mux2_1 _416_ (.A0(\scan_chain.scan_cells[20].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[19].scan_cell.data_out ),
    .S(net21),
    .X(_208_));
 sky130_fd_sc_hd__mux2_1 _417_ (.A0(\scan_chain.scan_cells[20].scan_cell.primary_ff ),
    .A1(_208_),
    .S(net34),
    .X(_128_));
 sky130_fd_sc_hd__mux2_1 _418_ (.A0(\dout[20] ),
    .A1(\scan_chain.scan_cells[20].scan_cell.primary_ff ),
    .S(net21),
    .X(_209_));
 sky130_fd_sc_hd__mux2_1 _419_ (.A0(\scan_chain.scan_cells[20].scan_cell.data_out ),
    .A1(_209_),
    .S(net35),
    .X(_129_));
 sky130_fd_sc_hd__mux2_1 _420_ (.A0(\scan_chain.scan_cells[1].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[0].scan_cell.data_out ),
    .S(net10),
    .X(_210_));
 sky130_fd_sc_hd__mux2_1 _421_ (.A0(\scan_chain.scan_cells[1].scan_cell.primary_ff ),
    .A1(_210_),
    .S(net23),
    .X(_130_));
 sky130_fd_sc_hd__mux2_1 _422_ (.A0(\dout[19] ),
    .A1(\scan_chain.scan_cells[19].scan_cell.primary_ff ),
    .S(net17),
    .X(_211_));
 sky130_fd_sc_hd__mux2_1 _423_ (.A0(\scan_chain.scan_cells[19].scan_cell.data_out ),
    .A1(_211_),
    .S(net32),
    .X(_131_));
 sky130_fd_sc_hd__mux2_1 _424_ (.A0(\scan_chain.scan_cells[18].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[17].scan_cell.data_out ),
    .S(net19),
    .X(_212_));
 sky130_fd_sc_hd__mux2_1 _425_ (.A0(\scan_chain.scan_cells[18].scan_cell.primary_ff ),
    .A1(_212_),
    .S(net31),
    .X(_132_));
 sky130_fd_sc_hd__mux2_1 _426_ (.A0(\dout[18] ),
    .A1(\scan_chain.scan_cells[18].scan_cell.primary_ff ),
    .S(net19),
    .X(_213_));
 sky130_fd_sc_hd__mux2_1 _427_ (.A0(\scan_chain.scan_cells[18].scan_cell.data_out ),
    .A1(_213_),
    .S(net31),
    .X(_133_));
 sky130_fd_sc_hd__mux2_1 _428_ (.A0(\scan_chain.scan_cells[17].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[16].scan_cell.data_out ),
    .S(net13),
    .X(_214_));
 sky130_fd_sc_hd__mux2_1 _429_ (.A0(\scan_chain.scan_cells[17].scan_cell.primary_ff ),
    .A1(_214_),
    .S(net31),
    .X(_134_));
 sky130_fd_sc_hd__mux2_1 _430_ (.A0(\dout[17] ),
    .A1(\scan_chain.scan_cells[17].scan_cell.primary_ff ),
    .S(net13),
    .X(_215_));
 sky130_fd_sc_hd__mux2_1 _431_ (.A0(\scan_chain.scan_cells[17].scan_cell.data_out ),
    .A1(_215_),
    .S(net31),
    .X(_135_));
 sky130_fd_sc_hd__mux2_1 _432_ (.A0(\scan_chain.scan_cells[16].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[15].scan_cell.data_out ),
    .S(net13),
    .X(_216_));
 sky130_fd_sc_hd__mux2_1 _433_ (.A0(\scan_chain.scan_cells[16].scan_cell.primary_ff ),
    .A1(_216_),
    .S(net28),
    .X(_136_));
 sky130_fd_sc_hd__mux2_1 _434_ (.A0(\dout[16] ),
    .A1(\scan_chain.scan_cells[16].scan_cell.primary_ff ),
    .S(net13),
    .X(_217_));
 sky130_fd_sc_hd__mux2_1 _435_ (.A0(\scan_chain.scan_cells[16].scan_cell.data_out ),
    .A1(_217_),
    .S(net28),
    .X(_137_));
 sky130_fd_sc_hd__mux2_1 _436_ (.A0(\scan_chain.scan_cells[15].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[14].scan_cell.data_out ),
    .S(net14),
    .X(_218_));
 sky130_fd_sc_hd__mux2_1 _437_ (.A0(\scan_chain.scan_cells[15].scan_cell.primary_ff ),
    .A1(_218_),
    .S(net28),
    .X(_138_));
 sky130_fd_sc_hd__mux2_1 _438_ (.A0(\dout[15] ),
    .A1(\scan_chain.scan_cells[15].scan_cell.primary_ff ),
    .S(net14),
    .X(_219_));
 sky130_fd_sc_hd__mux2_1 _439_ (.A0(\scan_chain.scan_cells[15].scan_cell.data_out ),
    .A1(_219_),
    .S(net28),
    .X(_139_));
 sky130_fd_sc_hd__mux2_1 _440_ (.A0(\scan_chain.scan_cells[14].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[13].scan_cell.data_out ),
    .S(net13),
    .X(_220_));
 sky130_fd_sc_hd__mux2_1 _441_ (.A0(\scan_chain.scan_cells[14].scan_cell.primary_ff ),
    .A1(_220_),
    .S(net28),
    .X(_140_));
 sky130_fd_sc_hd__mux2_1 _442_ (.A0(\dout[14] ),
    .A1(\scan_chain.scan_cells[14].scan_cell.primary_ff ),
    .S(net13),
    .X(_221_));
 sky130_fd_sc_hd__mux2_1 _443_ (.A0(\scan_chain.scan_cells[14].scan_cell.data_out ),
    .A1(_221_),
    .S(net28),
    .X(_141_));
 sky130_fd_sc_hd__mux2_1 _444_ (.A0(\scan_chain.scan_cells[13].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[12].scan_cell.data_out ),
    .S(net14),
    .X(_222_));
 sky130_fd_sc_hd__mux2_1 _445_ (.A0(\scan_chain.scan_cells[13].scan_cell.primary_ff ),
    .A1(_222_),
    .S(net28),
    .X(_142_));
 sky130_fd_sc_hd__mux2_1 _446_ (.A0(\dout[13] ),
    .A1(\scan_chain.scan_cells[13].scan_cell.primary_ff ),
    .S(net14),
    .X(_223_));
 sky130_fd_sc_hd__mux2_1 _447_ (.A0(\scan_chain.scan_cells[13].scan_cell.data_out ),
    .A1(_223_),
    .S(net28),
    .X(_143_));
 sky130_fd_sc_hd__mux2_1 _448_ (.A0(\scan_chain.scan_cells[12].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[11].scan_cell.data_out ),
    .S(net16),
    .X(_224_));
 sky130_fd_sc_hd__mux2_1 _449_ (.A0(\scan_chain.scan_cells[12].scan_cell.primary_ff ),
    .A1(_224_),
    .S(net30),
    .X(_000_));
 sky130_fd_sc_hd__mux2_1 _450_ (.A0(\dout[12] ),
    .A1(\scan_chain.scan_cells[12].scan_cell.primary_ff ),
    .S(net16),
    .X(_225_));
 sky130_fd_sc_hd__mux2_1 _451_ (.A0(\scan_chain.scan_cells[12].scan_cell.data_out ),
    .A1(_225_),
    .S(net37),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _452_ (.A0(\scan_chain.scan_cells[11].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[10].scan_cell.data_out ),
    .S(net16),
    .X(_226_));
 sky130_fd_sc_hd__mux2_1 _453_ (.A0(\scan_chain.scan_cells[11].scan_cell.primary_ff ),
    .A1(_226_),
    .S(net30),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _454_ (.A0(\dout[11] ),
    .A1(\scan_chain.scan_cells[11].scan_cell.primary_ff ),
    .S(net16),
    .X(_227_));
 sky130_fd_sc_hd__mux2_1 _455_ (.A0(\scan_chain.scan_cells[11].scan_cell.data_out ),
    .A1(_227_),
    .S(net30),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _456_ (.A0(\scan_chain.scan_cells[10].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[10].scan_cell.scan_in ),
    .S(net12),
    .X(_228_));
 sky130_fd_sc_hd__mux2_1 _457_ (.A0(\scan_chain.scan_cells[10].scan_cell.primary_ff ),
    .A1(_228_),
    .S(net29),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _458_ (.A0(\dout[10] ),
    .A1(\scan_chain.scan_cells[10].scan_cell.primary_ff ),
    .S(net13),
    .X(_229_));
 sky130_fd_sc_hd__mux2_1 _459_ (.A0(\scan_chain.scan_cells[10].scan_cell.data_out ),
    .A1(_229_),
    .S(net29),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _460_ (.A0(\scan_chain.scan_cells[0].scan_cell.data_out ),
    .A1(net2),
    .S(net10),
    .X(_230_));
 sky130_fd_sc_hd__mux2_1 _461_ (.A0(\scan_chain.scan_cells[0].scan_cell.primary_ff ),
    .A1(_230_),
    .S(net24),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _462_ (.A0(\dout[9] ),
    .A1(\scan_chain.scan_cells[9].scan_cell.primary_ff ),
    .S(net12),
    .X(_231_));
 sky130_fd_sc_hd__mux2_1 _463_ (.A0(\scan_chain.scan_cells[10].scan_cell.scan_in ),
    .A1(_231_),
    .S(net27),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _464_ (.A0(\scan_chain.scan_cells[8].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[7].scan_cell.data_out ),
    .S(net12),
    .X(_232_));
 sky130_fd_sc_hd__mux2_1 _465_ (.A0(\scan_chain.scan_cells[8].scan_cell.primary_ff ),
    .A1(_232_),
    .S(net27),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _466_ (.A0(\dout[8] ),
    .A1(\scan_chain.scan_cells[8].scan_cell.primary_ff ),
    .S(net15),
    .X(_233_));
 sky130_fd_sc_hd__mux2_1 _467_ (.A0(\scan_chain.scan_cells[8].scan_cell.data_out ),
    .A1(_233_),
    .S(net27),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _468_ (.A0(\scan_chain.scan_cells[7].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[6].scan_cell.data_out ),
    .S(net10),
    .X(_234_));
 sky130_fd_sc_hd__mux2_1 _469_ (.A0(\scan_chain.scan_cells[7].scan_cell.primary_ff ),
    .A1(_234_),
    .S(net29),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _470_ (.A0(\dout[7] ),
    .A1(\scan_chain.scan_cells[7].scan_cell.primary_ff ),
    .S(net15),
    .X(_235_));
 sky130_fd_sc_hd__mux2_1 _471_ (.A0(\scan_chain.scan_cells[7].scan_cell.data_out ),
    .A1(_235_),
    .S(net29),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _472_ (.A0(\scan_chain.scan_cells[71].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[70].scan_cell.data_in ),
    .S(net15),
    .X(_236_));
 sky130_fd_sc_hd__mux2_1 _473_ (.A0(\scan_chain.scan_cells[71].scan_cell.primary_ff ),
    .A1(_236_),
    .S(net25),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _474_ (.A0(\dout[6] ),
    .A1(\scan_chain.scan_cells[6].scan_cell.primary_ff ),
    .S(net11),
    .X(_237_));
 sky130_fd_sc_hd__mux2_1 _475_ (.A0(\scan_chain.scan_cells[6].scan_cell.data_out ),
    .A1(_237_),
    .S(net24),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _476_ (.A0(\scan_chain.scan_cells[69].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[68].scan_cell.data_in ),
    .S(net15),
    .X(_238_));
 sky130_fd_sc_hd__mux2_1 _477_ (.A0(\scan_chain.scan_cells[69].scan_cell.primary_ff ),
    .A1(_238_),
    .S(net25),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _478_ (.A0(\dout[5] ),
    .A1(\scan_chain.scan_cells[5].scan_cell.primary_ff ),
    .S(net11),
    .X(_239_));
 sky130_fd_sc_hd__mux2_1 _479_ (.A0(\scan_chain.scan_cells[5].scan_cell.data_out ),
    .A1(_239_),
    .S(net24),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _480_ (.A0(\scan_chain.scan_cells[59].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[58].scan_cell.data_in ),
    .S(net19),
    .X(_240_));
 sky130_fd_sc_hd__mux2_1 _481_ (.A0(\scan_chain.scan_cells[59].scan_cell.primary_ff ),
    .A1(_240_),
    .S(net36),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _482_ (.A0(\dout[4] ),
    .A1(\scan_chain.scan_cells[4].scan_cell.primary_ff ),
    .S(net10),
    .X(_241_));
 sky130_fd_sc_hd__mux2_1 _483_ (.A0(\scan_chain.scan_cells[4].scan_cell.data_out ),
    .A1(_241_),
    .S(net23),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _484_ (.A0(\scan_chain.scan_cells[49].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[48].scan_cell.data_in ),
    .S(net17),
    .X(_242_));
 sky130_fd_sc_hd__mux2_1 _485_ (.A0(\scan_chain.scan_cells[49].scan_cell.primary_ff ),
    .A1(_242_),
    .S(net31),
    .X(_018_));
 sky130_fd_sc_hd__mux2_1 _486_ (.A0(\dout[3] ),
    .A1(\scan_chain.scan_cells[3].scan_cell.primary_ff ),
    .S(net10),
    .X(_243_));
 sky130_fd_sc_hd__mux2_1 _487_ (.A0(\scan_chain.scan_cells[3].scan_cell.data_out ),
    .A1(_243_),
    .S(net23),
    .X(_019_));
 sky130_fd_sc_hd__mux2_1 _488_ (.A0(\scan_chain.scan_cells[39].scan_cell.data_in ),
    .A1(\scan_chain.scan_cells[38].scan_cell.data_in ),
    .S(net11),
    .X(_244_));
 sky130_fd_sc_hd__mux2_1 _489_ (.A0(\scan_chain.scan_cells[39].scan_cell.primary_ff ),
    .A1(_244_),
    .S(net24),
    .X(_020_));
 sky130_fd_sc_hd__mux2_1 _490_ (.A0(\dout[2] ),
    .A1(\scan_chain.scan_cells[2].scan_cell.primary_ff ),
    .S(net10),
    .X(_245_));
 sky130_fd_sc_hd__mux2_1 _491_ (.A0(\scan_chain.scan_cells[2].scan_cell.data_out ),
    .A1(_245_),
    .S(net23),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _492_ (.A0(\scan_chain.scan_cells[29].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[28].scan_cell.data_out ),
    .S(net18),
    .X(_246_));
 sky130_fd_sc_hd__mux2_1 _493_ (.A0(\scan_chain.scan_cells[29].scan_cell.primary_ff ),
    .A1(_246_),
    .S(net33),
    .X(_022_));
 sky130_fd_sc_hd__mux2_1 _494_ (.A0(\dout[1] ),
    .A1(\scan_chain.scan_cells[1].scan_cell.primary_ff ),
    .S(net10),
    .X(_247_));
 sky130_fd_sc_hd__mux2_1 _495_ (.A0(\scan_chain.scan_cells[1].scan_cell.data_out ),
    .A1(_247_),
    .S(net23),
    .X(_023_));
 sky130_fd_sc_hd__mux2_1 _496_ (.A0(\scan_chain.scan_cells[19].scan_cell.data_out ),
    .A1(\scan_chain.scan_cells[18].scan_cell.data_out ),
    .S(net19),
    .X(_248_));
 sky130_fd_sc_hd__mux2_1 _497_ (.A0(\scan_chain.scan_cells[19].scan_cell.primary_ff ),
    .A1(_248_),
    .S(net31),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _498_ (.A0(\dout[0] ),
    .A1(\scan_chain.scan_cells[0].scan_cell.primary_ff ),
    .S(net11),
    .X(_249_));
 sky130_fd_sc_hd__mux2_1 _499_ (.A0(\scan_chain.scan_cells[0].scan_cell.data_out ),
    .A1(_249_),
    .S(net24),
    .X(_025_));
 sky130_fd_sc_hd__dfrtp_1 _500_ (.CLK(clknet_3_0__leaf_ui_in[3]),
    .D(_026_),
    .RESET_B(net43),
    .Q(\scan_chain.scan_cells[9].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _501_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_027_),
    .RESET_B(net38),
    .Q(\scan_chain.scan_cells[71].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _502_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_028_),
    .RESET_B(net38),
    .Q(\scan_chain.scan_cells[70].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _503_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_029_),
    .RESET_B(net38),
    .Q(\scan_chain.scan_cells[70].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _504_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_030_),
    .RESET_B(net43),
    .Q(\scan_chain.scan_cells[6].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _505_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_031_),
    .RESET_B(net38),
    .Q(\scan_chain.scan_cells[69].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _506_ (.CLK(clknet_3_2__leaf_ui_in[3]),
    .D(_032_),
    .RESET_B(net39),
    .Q(\scan_chain.scan_cells[68].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _507_ (.CLK(clknet_3_2__leaf_ui_in[4]),
    .D(_033_),
    .RESET_B(net39),
    .Q(\scan_chain.scan_cells[68].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _508_ (.CLK(clknet_3_2__leaf_ui_in[3]),
    .D(_034_),
    .RESET_B(net39),
    .Q(\scan_chain.scan_cells[67].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _509_ (.CLK(clknet_3_2__leaf_ui_in[4]),
    .D(_035_),
    .RESET_B(net39),
    .Q(\scan_chain.scan_cells[67].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _510_ (.CLK(clknet_3_2__leaf_ui_in[3]),
    .D(_036_),
    .RESET_B(net39),
    .Q(\scan_chain.scan_cells[66].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _511_ (.CLK(clknet_3_2__leaf_ui_in[4]),
    .D(_037_),
    .RESET_B(net39),
    .Q(\scan_chain.scan_cells[66].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _512_ (.CLK(clknet_3_7__leaf_ui_in[3]),
    .D(_038_),
    .RESET_B(net54),
    .Q(\scan_chain.scan_cells[65].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _513_ (.CLK(clknet_3_4__leaf_ui_in[4]),
    .D(_039_),
    .RESET_B(net54),
    .Q(\scan_chain.scan_cells[65].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _514_ (.CLK(clknet_3_7__leaf_ui_in[3]),
    .D(_040_),
    .RESET_B(net54),
    .Q(\scan_chain.scan_cells[64].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _515_ (.CLK(clknet_3_4__leaf_ui_in[4]),
    .D(_041_),
    .RESET_B(net54),
    .Q(\scan_chain.scan_cells[64].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _516_ (.CLK(clknet_3_4__leaf_ui_in[3]),
    .D(_042_),
    .RESET_B(net53),
    .Q(\scan_chain.scan_cells[63].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _517_ (.CLK(clknet_3_4__leaf_ui_in[4]),
    .D(_043_),
    .RESET_B(net53),
    .Q(\scan_chain.scan_cells[63].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _518_ (.CLK(clknet_3_4__leaf_ui_in[3]),
    .D(_044_),
    .RESET_B(net53),
    .Q(\scan_chain.scan_cells[62].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _519_ (.CLK(clknet_3_4__leaf_ui_in[4]),
    .D(_045_),
    .RESET_B(net53),
    .Q(\scan_chain.scan_cells[62].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _520_ (.CLK(clknet_3_4__leaf_ui_in[3]),
    .D(_046_),
    .RESET_B(net53),
    .Q(\scan_chain.scan_cells[61].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _521_ (.CLK(clknet_3_4__leaf_ui_in[4]),
    .D(_047_),
    .RESET_B(net53),
    .Q(\scan_chain.scan_cells[61].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _522_ (.CLK(clknet_3_7__leaf_ui_in[3]),
    .D(_048_),
    .RESET_B(net53),
    .Q(\scan_chain.scan_cells[60].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _523_ (.CLK(clknet_3_7__leaf_ui_in[4]),
    .D(_049_),
    .RESET_B(net53),
    .Q(\scan_chain.scan_cells[60].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _524_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_050_),
    .RESET_B(net40),
    .Q(\scan_chain.scan_cells[5].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _525_ (.CLK(clknet_3_7__leaf_ui_in[4]),
    .D(_051_),
    .RESET_B(net54),
    .Q(\scan_chain.scan_cells[59].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _526_ (.CLK(clknet_3_7__leaf_ui_in[3]),
    .D(_052_),
    .RESET_B(net54),
    .Q(\scan_chain.scan_cells[58].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _527_ (.CLK(clknet_3_7__leaf_ui_in[4]),
    .D(_053_),
    .RESET_B(net54),
    .Q(\scan_chain.scan_cells[58].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _528_ (.CLK(clknet_3_7__leaf_ui_in[3]),
    .D(_054_),
    .RESET_B(net51),
    .Q(\scan_chain.scan_cells[57].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _529_ (.CLK(clknet_3_7__leaf_ui_in[4]),
    .D(_055_),
    .RESET_B(net51),
    .Q(\scan_chain.scan_cells[57].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _530_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_056_),
    .RESET_B(net52),
    .Q(\scan_chain.scan_cells[56].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _531_ (.CLK(clknet_3_7__leaf_ui_in[4]),
    .D(_057_),
    .RESET_B(net52),
    .Q(\scan_chain.scan_cells[56].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _532_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_058_),
    .RESET_B(net51),
    .Q(\scan_chain.scan_cells[55].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_2 _533_ (.CLK(clknet_3_7__leaf_ui_in[4]),
    .D(_059_),
    .RESET_B(net51),
    .Q(\scan_chain.scan_cells[55].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _534_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_060_),
    .RESET_B(net51),
    .Q(\scan_chain.scan_cells[54].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_2 _535_ (.CLK(clknet_3_7__leaf_ui_in[4]),
    .D(_061_),
    .RESET_B(net51),
    .Q(\scan_chain.scan_cells[54].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _536_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_062_),
    .RESET_B(net51),
    .Q(\scan_chain.scan_cells[53].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_2 _537_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_063_),
    .RESET_B(net51),
    .Q(\scan_chain.scan_cells[53].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _538_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_064_),
    .RESET_B(net50),
    .Q(\scan_chain.scan_cells[52].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_2 _539_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_065_),
    .RESET_B(net52),
    .Q(\scan_chain.scan_cells[52].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _540_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_066_),
    .RESET_B(net48),
    .Q(\scan_chain.scan_cells[51].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_2 _541_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_067_),
    .RESET_B(net48),
    .Q(\scan_chain.scan_cells[51].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _542_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_068_),
    .RESET_B(net48),
    .Q(\scan_chain.scan_cells[50].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _543_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_069_),
    .RESET_B(net49),
    .Q(\scan_chain.scan_cells[50].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _544_ (.CLK(clknet_3_2__leaf_ui_in[3]),
    .D(_070_),
    .RESET_B(net40),
    .Q(\scan_chain.scan_cells[4].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _545_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_071_),
    .RESET_B(net50),
    .Q(\scan_chain.scan_cells[49].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _546_ (.CLK(clknet_3_1__leaf_ui_in[3]),
    .D(_072_),
    .RESET_B(net48),
    .Q(\scan_chain.scan_cells[48].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _547_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_073_),
    .RESET_B(net48),
    .Q(\scan_chain.scan_cells[48].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _548_ (.CLK(clknet_3_1__leaf_ui_in[3]),
    .D(_074_),
    .RESET_B(net45),
    .Q(\scan_chain.scan_cells[47].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _549_ (.CLK(clknet_3_1__leaf_ui_in[4]),
    .D(_075_),
    .RESET_B(net45),
    .Q(\scan_chain.scan_cells[47].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _550_ (.CLK(clknet_3_0__leaf_ui_in[3]),
    .D(_076_),
    .RESET_B(net45),
    .Q(\scan_chain.scan_cells[46].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _551_ (.CLK(clknet_3_1__leaf_ui_in[4]),
    .D(_077_),
    .RESET_B(net45),
    .Q(\scan_chain.scan_cells[46].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _552_ (.CLK(clknet_3_0__leaf_ui_in[3]),
    .D(_078_),
    .RESET_B(net43),
    .Q(\scan_chain.scan_cells[45].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _553_ (.CLK(clknet_3_0__leaf_ui_in[4]),
    .D(_079_),
    .RESET_B(net45),
    .Q(\scan_chain.scan_cells[45].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _554_ (.CLK(clknet_3_0__leaf_ui_in[3]),
    .D(_080_),
    .RESET_B(net46),
    .Q(\scan_chain.scan_cells[44].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _555_ (.CLK(clknet_3_1__leaf_ui_in[4]),
    .D(_081_),
    .RESET_B(net46),
    .Q(\scan_chain.scan_cells[44].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _556_ (.CLK(clknet_3_0__leaf_ui_in[3]),
    .D(_082_),
    .RESET_B(net43),
    .Q(\scan_chain.scan_cells[43].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _557_ (.CLK(clknet_3_0__leaf_ui_in[4]),
    .D(_083_),
    .RESET_B(net44),
    .Q(\scan_chain.scan_cells[43].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _558_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_084_),
    .RESET_B(net44),
    .Q(\scan_chain.scan_cells[42].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _559_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_085_),
    .RESET_B(net44),
    .Q(\scan_chain.scan_cells[42].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _560_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_086_),
    .RESET_B(net43),
    .Q(\scan_chain.scan_cells[41].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _561_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_087_),
    .RESET_B(net43),
    .Q(\scan_chain.scan_cells[41].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _562_ (.CLK(clknet_3_0__leaf_ui_in[3]),
    .D(_088_),
    .RESET_B(net43),
    .Q(\scan_chain.scan_cells[40].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _563_ (.CLK(clknet_3_0__leaf_ui_in[4]),
    .D(_089_),
    .RESET_B(net44),
    .Q(\scan_chain.scan_cells[40].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _564_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_090_),
    .RESET_B(net40),
    .Q(\scan_chain.scan_cells[3].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _565_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_091_),
    .RESET_B(net40),
    .Q(\scan_chain.scan_cells[39].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _566_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_092_),
    .RESET_B(net42),
    .Q(\scan_chain.scan_cells[38].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _567_ (.CLK(clknet_3_2__leaf_ui_in[4]),
    .D(_093_),
    .RESET_B(net42),
    .Q(\scan_chain.scan_cells[38].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _568_ (.CLK(clknet_3_2__leaf_ui_in[3]),
    .D(_094_),
    .RESET_B(net42),
    .Q(\scan_chain.scan_cells[37].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _569_ (.CLK(clknet_3_2__leaf_ui_in[4]),
    .D(_095_),
    .RESET_B(net42),
    .Q(\scan_chain.scan_cells[37].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _570_ (.CLK(clknet_3_2__leaf_ui_in[3]),
    .D(_096_),
    .RESET_B(net40),
    .Q(\scan_chain.scan_cells[36].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _571_ (.CLK(clknet_3_2__leaf_ui_in[4]),
    .D(_097_),
    .RESET_B(net42),
    .Q(\scan_chain.scan_cells[36].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _572_ (.CLK(clknet_3_2__leaf_ui_in[3]),
    .D(_098_),
    .RESET_B(net38),
    .Q(\scan_chain.scan_cells[35].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_2 _573_ (.CLK(clknet_3_2__leaf_ui_in[4]),
    .D(_099_),
    .RESET_B(net38),
    .Q(\scan_chain.scan_cells[35].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _574_ (.CLK(clknet_3_2__leaf_ui_in[3]),
    .D(_100_),
    .RESET_B(net38),
    .Q(\scan_chain.scan_cells[34].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_2 _575_ (.CLK(clknet_3_2__leaf_ui_in[4]),
    .D(_101_),
    .RESET_B(net38),
    .Q(\scan_chain.scan_cells[34].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _576_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_102_),
    .RESET_B(net39),
    .Q(\scan_chain.scan_cells[33].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_2 _577_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_103_),
    .RESET_B(net39),
    .Q(\scan_chain.scan_cells[33].scan_cell.data_in ));
 sky130_fd_sc_hd__dfrtp_1 _578_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_104_),
    .RESET_B(net49),
    .Q(\scan_chain.scan_cells[32].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _579_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_105_),
    .RESET_B(net49),
    .Q(\scan_chain.scan_cells[32].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _580_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_106_),
    .RESET_B(net49),
    .Q(\scan_chain.scan_cells[31].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _581_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_107_),
    .RESET_B(net49),
    .Q(\scan_chain.scan_cells[31].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _582_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_108_),
    .RESET_B(net51),
    .Q(\scan_chain.scan_cells[30].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _583_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_109_),
    .RESET_B(net51),
    .Q(\scan_chain.scan_cells[30].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _584_ (.CLK(clknet_3_2__leaf_ui_in[3]),
    .D(_110_),
    .RESET_B(net40),
    .Q(\scan_chain.scan_cells[2].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _585_ (.CLK(clknet_3_7__leaf_ui_in[4]),
    .D(_111_),
    .RESET_B(net52),
    .Q(\scan_chain.scan_cells[29].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _586_ (.CLK(clknet_3_4__leaf_ui_in[3]),
    .D(_112_),
    .RESET_B(net53),
    .Q(\scan_chain.scan_cells[28].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _587_ (.CLK(clknet_3_7__leaf_ui_in[4]),
    .D(_113_),
    .RESET_B(net53),
    .Q(\scan_chain.scan_cells[28].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _588_ (.CLK(clknet_3_4__leaf_ui_in[3]),
    .D(_114_),
    .RESET_B(net54),
    .Q(\scan_chain.scan_cells[27].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _589_ (.CLK(clknet_3_4__leaf_ui_in[4]),
    .D(_115_),
    .RESET_B(net54),
    .Q(\scan_chain.scan_cells[27].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _590_ (.CLK(clknet_3_5__leaf_ui_in[3]),
    .D(_116_),
    .RESET_B(net47),
    .Q(\scan_chain.scan_cells[26].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _591_ (.CLK(clknet_3_5__leaf_ui_in[4]),
    .D(_117_),
    .RESET_B(net47),
    .Q(\scan_chain.scan_cells[26].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _592_ (.CLK(clknet_3_5__leaf_ui_in[3]),
    .D(_118_),
    .RESET_B(net47),
    .Q(\scan_chain.scan_cells[25].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _593_ (.CLK(clknet_3_5__leaf_ui_in[4]),
    .D(_119_),
    .RESET_B(net47),
    .Q(\scan_chain.scan_cells[25].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _594_ (.CLK(clknet_3_5__leaf_ui_in[3]),
    .D(_120_),
    .RESET_B(net47),
    .Q(\scan_chain.scan_cells[24].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _595_ (.CLK(clknet_3_5__leaf_ui_in[4]),
    .D(_121_),
    .RESET_B(net47),
    .Q(\scan_chain.scan_cells[24].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _596_ (.CLK(clknet_3_5__leaf_ui_in[3]),
    .D(_122_),
    .RESET_B(net47),
    .Q(\scan_chain.scan_cells[23].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _597_ (.CLK(clknet_3_5__leaf_ui_in[4]),
    .D(_123_),
    .RESET_B(net56),
    .Q(\scan_chain.scan_cells[23].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _598_ (.CLK(clknet_3_5__leaf_ui_in[3]),
    .D(_124_),
    .RESET_B(net55),
    .Q(\scan_chain.scan_cells[22].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _599_ (.CLK(clknet_3_5__leaf_ui_in[4]),
    .D(_125_),
    .RESET_B(net55),
    .Q(\scan_chain.scan_cells[22].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _600_ (.CLK(clknet_3_4__leaf_ui_in[3]),
    .D(_126_),
    .RESET_B(net55),
    .Q(\scan_chain.scan_cells[21].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _601_ (.CLK(clknet_3_4__leaf_ui_in[4]),
    .D(_127_),
    .RESET_B(net55),
    .Q(\scan_chain.scan_cells[21].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _602_ (.CLK(clknet_3_7__leaf_ui_in[3]),
    .D(_128_),
    .RESET_B(net55),
    .Q(\scan_chain.scan_cells[20].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _603_ (.CLK(clknet_3_4__leaf_ui_in[4]),
    .D(_129_),
    .RESET_B(net55),
    .Q(\scan_chain.scan_cells[20].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _604_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_130_),
    .RESET_B(net41),
    .Q(\scan_chain.scan_cells[1].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _605_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_131_),
    .RESET_B(net50),
    .Q(\scan_chain.scan_cells[19].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _606_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_132_),
    .RESET_B(net48),
    .Q(\scan_chain.scan_cells[18].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _607_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_133_),
    .RESET_B(net48),
    .Q(\scan_chain.scan_cells[18].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _608_ (.CLK(clknet_3_1__leaf_ui_in[3]),
    .D(_134_),
    .RESET_B(net48),
    .Q(\scan_chain.scan_cells[17].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _609_ (.CLK(clknet_3_6__leaf_ui_in[4]),
    .D(_135_),
    .RESET_B(net48),
    .Q(\scan_chain.scan_cells[17].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _610_ (.CLK(clknet_3_1__leaf_ui_in[3]),
    .D(_136_),
    .RESET_B(net45),
    .Q(\scan_chain.scan_cells[16].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _611_ (.CLK(clknet_3_1__leaf_ui_in[4]),
    .D(_137_),
    .RESET_B(net45),
    .Q(\scan_chain.scan_cells[16].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _612_ (.CLK(clknet_3_1__leaf_ui_in[3]),
    .D(_138_),
    .RESET_B(net45),
    .Q(\scan_chain.scan_cells[15].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _613_ (.CLK(clknet_3_1__leaf_ui_in[4]),
    .D(_139_),
    .RESET_B(net46),
    .Q(\scan_chain.scan_cells[15].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _614_ (.CLK(clknet_3_1__leaf_ui_in[3]),
    .D(_140_),
    .RESET_B(net46),
    .Q(\scan_chain.scan_cells[14].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _615_ (.CLK(clknet_3_1__leaf_ui_in[4]),
    .D(_141_),
    .RESET_B(net46),
    .Q(\scan_chain.scan_cells[14].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _616_ (.CLK(clknet_3_1__leaf_ui_in[3]),
    .D(_142_),
    .RESET_B(net46),
    .Q(\scan_chain.scan_cells[13].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _617_ (.CLK(clknet_3_1__leaf_ui_in[4]),
    .D(_143_),
    .RESET_B(net46),
    .Q(\scan_chain.scan_cells[13].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _618_ (.CLK(clknet_3_5__leaf_ui_in[3]),
    .D(_000_),
    .RESET_B(net47),
    .Q(\scan_chain.scan_cells[12].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _619_ (.CLK(clknet_3_5__leaf_ui_in[4]),
    .D(_001_),
    .RESET_B(net56),
    .Q(\scan_chain.scan_cells[12].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _620_ (.CLK(clknet_3_5__leaf_ui_in[3]),
    .D(_002_),
    .RESET_B(net47),
    .Q(\scan_chain.scan_cells[11].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _621_ (.CLK(clknet_3_5__leaf_ui_in[4]),
    .D(_003_),
    .RESET_B(net47),
    .Q(\scan_chain.scan_cells[11].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _622_ (.CLK(clknet_3_0__leaf_ui_in[3]),
    .D(_004_),
    .RESET_B(net45),
    .Q(\scan_chain.scan_cells[10].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_4 _623_ (.CLK(clknet_3_1__leaf_ui_in[4]),
    .D(_005_),
    .RESET_B(net45),
    .Q(\scan_chain.scan_cells[10].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _624_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_006_),
    .RESET_B(net41),
    .Q(\scan_chain.scan_cells[0].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _625_ (.CLK(clknet_3_0__leaf_ui_in[4]),
    .D(_007_),
    .RESET_B(net44),
    .Q(\scan_chain.scan_cells[10].scan_cell.scan_in ));
 sky130_fd_sc_hd__dfrtp_1 _626_ (.CLK(clknet_3_0__leaf_ui_in[3]),
    .D(_008_),
    .RESET_B(net44),
    .Q(\scan_chain.scan_cells[8].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _627_ (.CLK(clknet_3_0__leaf_ui_in[4]),
    .D(_009_),
    .RESET_B(net44),
    .Q(\scan_chain.scan_cells[8].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _628_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_010_),
    .RESET_B(net43),
    .Q(\scan_chain.scan_cells[7].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _629_ (.CLK(clknet_3_0__leaf_ui_in[4]),
    .D(_011_),
    .RESET_B(net43),
    .Q(\scan_chain.scan_cells[7].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _630_ (.CLK(clknet_3_2__leaf_ui_in[3]),
    .D(_012_),
    .RESET_B(net38),
    .Q(\scan_chain.scan_cells[71].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _631_ (.CLK(clknet_3_0__leaf_ui_in[4]),
    .D(_013_),
    .RESET_B(net43),
    .Q(\scan_chain.scan_cells[6].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _632_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_014_),
    .RESET_B(net38),
    .Q(\scan_chain.scan_cells[69].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _633_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_015_),
    .RESET_B(net41),
    .Q(\scan_chain.scan_cells[5].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _634_ (.CLK(clknet_3_7__leaf_ui_in[3]),
    .D(_016_),
    .RESET_B(net52),
    .Q(\scan_chain.scan_cells[59].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _635_ (.CLK(clknet_3_2__leaf_ui_in[4]),
    .D(_017_),
    .RESET_B(net40),
    .Q(\scan_chain.scan_cells[4].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _636_ (.CLK(clknet_3_6__leaf_ui_in[3]),
    .D(_018_),
    .RESET_B(net48),
    .Q(\scan_chain.scan_cells[49].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _637_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_019_),
    .RESET_B(net40),
    .Q(\scan_chain.scan_cells[3].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _638_ (.CLK(clknet_3_3__leaf_ui_in[3]),
    .D(_020_),
    .RESET_B(net41),
    .Q(\scan_chain.scan_cells[39].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _639_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_021_),
    .RESET_B(net40),
    .Q(\scan_chain.scan_cells[2].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _640_ (.CLK(clknet_3_7__leaf_ui_in[3]),
    .D(_022_),
    .RESET_B(net52),
    .Q(\scan_chain.scan_cells[29].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _641_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_023_),
    .RESET_B(net40),
    .Q(\scan_chain.scan_cells[1].scan_cell.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _642_ (.CLK(clknet_3_1__leaf_ui_in[3]),
    .D(_024_),
    .RESET_B(net50),
    .Q(\scan_chain.scan_cells[19].scan_cell.primary_ff ));
 sky130_fd_sc_hd__dfrtp_1 _643_ (.CLK(clknet_3_3__leaf_ui_in[4]),
    .D(_025_),
    .RESET_B(net41),
    .Q(\scan_chain.scan_cells[0].scan_cell.data_out ));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_79 (.LO(net79));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_ui_in[3]  (.A(ui_in[3]),
    .X(clknet_0_ui_in[3]));
 sky130_fd_sc_hd__clkbuf_4 _666_ (.A(\scan_chain.scan_cells[71].scan_cell.data_in ),
    .X(uo_out[0]));
 sky130_fd_sc_hd__buf_2 _667_ (.A(\scan_chain.scan_cells[0].scan_cell.data_out ),
    .X(uo_out[1]));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_2_Left_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_2_Left_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_2_Left_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_2_Left_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_2_Left_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_2_Left_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_2_Left_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_2_Left_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_2_Left_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Left_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Left_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Left_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Left_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Left_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Left_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Left_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Left_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Left_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Left_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Left_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Left_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Left_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Left_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Left_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Left_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Left_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Left_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Left_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Left_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Left_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Left_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_2_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_2_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_2_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_2_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_2_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_2_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_2_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_2_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_2_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_2_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_2_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_361 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(rst_n),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 fanout5 (.A(net6),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 fanout6 (.A(_145_),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 fanout7 (.A(net8),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 fanout8 (.A(_145_),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 fanout9 (.A(net15),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 fanout10 (.A(net11),
    .X(net10));
 sky130_fd_sc_hd__buf_2 fanout11 (.A(net15),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 fanout12 (.A(net15),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 fanout13 (.A(net14),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 fanout14 (.A(net15),
    .X(net14));
 sky130_fd_sc_hd__buf_2 fanout15 (.A(net4),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 fanout16 (.A(net22),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 fanout17 (.A(net19),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 fanout18 (.A(net19),
    .X(net18));
 sky130_fd_sc_hd__buf_2 fanout19 (.A(net22),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 fanout20 (.A(net22),
    .X(net20));
 sky130_fd_sc_hd__buf_2 fanout21 (.A(net22),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 fanout22 (.A(net4),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 fanout23 (.A(net26),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 fanout24 (.A(net26),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 fanout25 (.A(net26),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 fanout26 (.A(net37),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 fanout27 (.A(net29),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 fanout28 (.A(net29),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 fanout29 (.A(net37),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 fanout30 (.A(net37),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 fanout31 (.A(net32),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 fanout32 (.A(net36),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 fanout33 (.A(net36),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 fanout34 (.A(net35),
    .X(net34));
 sky130_fd_sc_hd__buf_2 fanout35 (.A(net36),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 fanout36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 fanout37 (.A(net3),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_4 fanout38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__buf_2 fanout39 (.A(net57),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_4 fanout40 (.A(net42),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 fanout41 (.A(net42),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 fanout42 (.A(net57),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 fanout43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__buf_2 fanout44 (.A(net57),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 fanout45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__buf_2 fanout46 (.A(net57),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 fanout47 (.A(net56),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 fanout48 (.A(net50),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 fanout49 (.A(net50),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 fanout50 (.A(net56),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 fanout51 (.A(net52),
    .X(net51));
 sky130_fd_sc_hd__buf_2 fanout52 (.A(net56),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 fanout53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 fanout54 (.A(net55),
    .X(net54));
 sky130_fd_sc_hd__buf_2 fanout55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_4 fanout56 (.A(net57),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 fanout57 (.A(net1),
    .X(net57));
 sky130_fd_sc_hd__conb_1 tt_um_openram_top_58 (.LO(net58));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_0__f_ui_in[3]  (.A(clknet_0_ui_in[3]),
    .X(clknet_3_0__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_1__f_ui_in[3]  (.A(clknet_0_ui_in[3]),
    .X(clknet_3_1__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_2__f_ui_in[3]  (.A(clknet_0_ui_in[3]),
    .X(clknet_3_2__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_3__f_ui_in[3]  (.A(clknet_0_ui_in[3]),
    .X(clknet_3_3__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_4__f_ui_in[3]  (.A(clknet_0_ui_in[3]),
    .X(clknet_3_4__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_5__f_ui_in[3]  (.A(clknet_0_ui_in[3]),
    .X(clknet_3_5__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_6__f_ui_in[3]  (.A(clknet_0_ui_in[3]),
    .X(clknet_3_6__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_7__f_ui_in[3]  (.A(clknet_0_ui_in[3]),
    .X(clknet_3_7__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkinvlp_4 clkload0 (.A(clknet_3_0__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkinvlp_4 clkload1 (.A(clknet_3_1__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkinv_2 clkload2 (.A(clknet_3_2__leaf_ui_in[3]));
 sky130_fd_sc_hd__inv_6 clkload3 (.A(clknet_3_4__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkinv_4 clkload4 (.A(clknet_3_5__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkbuf_4 clkload5 (.A(clknet_3_6__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkinvlp_4 clkload6 (.A(clknet_3_7__leaf_ui_in[3]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_ui_in[4]  (.A(ui_in[4]),
    .X(clknet_0_ui_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_0__f_ui_in[4]  (.A(clknet_0_ui_in[4]),
    .X(clknet_3_0__leaf_ui_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_1__f_ui_in[4]  (.A(clknet_0_ui_in[4]),
    .X(clknet_3_1__leaf_ui_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_2__f_ui_in[4]  (.A(clknet_0_ui_in[4]),
    .X(clknet_3_2__leaf_ui_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_3__f_ui_in[4]  (.A(clknet_0_ui_in[4]),
    .X(clknet_3_3__leaf_ui_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_4__f_ui_in[4]  (.A(clknet_0_ui_in[4]),
    .X(clknet_3_4__leaf_ui_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_5__f_ui_in[4]  (.A(clknet_0_ui_in[4]),
    .X(clknet_3_5__leaf_ui_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_6__f_ui_in[4]  (.A(clknet_0_ui_in[4]),
    .X(clknet_3_6__leaf_ui_in[4]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_7__f_ui_in[4]  (.A(clknet_0_ui_in[4]),
    .X(clknet_3_7__leaf_ui_in[4]));
 sky130_fd_sc_hd__clkinvlp_4 clkload7 (.A(clknet_3_0__leaf_ui_in[4]));
 sky130_fd_sc_hd__bufinv_16 clkload8 (.A(clknet_3_1__leaf_ui_in[4]));
 sky130_fd_sc_hd__clkinv_2 clkload9 (.A(clknet_3_2__leaf_ui_in[4]));
 sky130_fd_sc_hd__clkbuf_4 clkload10 (.A(clknet_3_3__leaf_ui_in[4]));
 sky130_fd_sc_hd__bufinv_16 clkload11 (.A(clknet_3_4__leaf_ui_in[4]));
 sky130_fd_sc_hd__clkinvlp_4 clkload12 (.A(clknet_3_5__leaf_ui_in[4]));
 sky130_fd_sc_hd__clkinv_2 clkload13 (.A(clknet_3_7__leaf_ui_in[4]));
 assign uio_oe[0] = net58;
 assign uio_oe[1] = net59;
 assign uio_oe[2] = net60;
 assign uio_oe[3] = net61;
 assign uio_oe[4] = net62;
 assign uio_oe[5] = net63;
 assign uio_oe[6] = net64;
 assign uio_oe[7] = net65;
 assign uio_out[0] = net66;
 assign uio_out[1] = net67;
 assign uio_out[2] = net68;
 assign uio_out[3] = net69;
 assign uio_out[4] = net70;
 assign uio_out[5] = net71;
 assign uio_out[6] = net72;
 assign uio_out[7] = net73;
 assign uo_out[2] = net74;
 assign uo_out[3] = net75;
 assign uo_out[4] = net76;
 assign uo_out[5] = net77;
 assign uo_out[6] = net78;
 assign uo_out[7] = net79;
endmodule
